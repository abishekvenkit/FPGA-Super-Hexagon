module hsl_to_rgb(  input  logic Clk,
                    input  logic [5:0] Hue,
                    input  logic [3:0] Saturation,
                    input  logic [3:0] Luminance,
                    output logic [7:0] Red,
                    output logic [7:0] Green,
                    output logic [7:0] Blue
                    );

    reg signed [23:0] rgb [0:16383];
    logic [13:0] index;
    assign index = {Hue, Saturation, Luminance};
	 logic [23:0] rgb_val;

    always_ff @ (posedge Clk) begin
	     rgb_val <= rgb[index];
    end
	 
	 always_comb begin
	     Red = rgb_val[23:16];
		  Green = rgb_val[15:8];
		  Blue = rgb_val[7:0];
	 end

    initial begin
rgb[0] = 24'b000000000000000000000000;
rgb[1] = 24'b000100010001000100010001;
rgb[2] = 24'b001000100010001000100010;
rgb[3] = 24'b001100110011001100110011;
rgb[4] = 24'b010001000100010001000100;
rgb[5] = 24'b010101010101010101010101;
rgb[6] = 24'b011001100110011001100110;
rgb[7] = 24'b011101110111011101110111;
rgb[8] = 24'b100010001000100010001000;
rgb[9] = 24'b100110011001100110011001;
rgb[10] = 24'b101010101010101010101010;
rgb[11] = 24'b101110111011101110111011;
rgb[12] = 24'b110011001100110011001100;
rgb[13] = 24'b110111011101110111011101;
rgb[14] = 24'b111011101110111011101110;
rgb[15] = 24'b111111111111111111111111;
rgb[16] = 24'b000000000000000000000000;
rgb[17] = 24'b000100100000111100001111;
rgb[18] = 24'b001001000001111100011111;
rgb[19] = 24'b001101100010111100101111;
rgb[20] = 24'b010010000011111100111111;
rgb[21] = 24'b010110100100111101001111;
rgb[22] = 24'b011011000101111101011111;
rgb[23] = 24'b011111100110111101101111;
rgb[24] = 24'b100011111000000010000000;
rgb[25] = 24'b100111111001001010010010;
rgb[26] = 24'b101011111010010010100100;
rgb[27] = 24'b101111111011011010110110;
rgb[28] = 24'b110011111100100011001000;
rgb[29] = 24'b110111111101101011011010;
rgb[30] = 24'b111011111110110011101100;
rgb[31] = 24'b111111111111111111111111;
rgb[32] = 24'b000000000000000000000000;
rgb[33] = 24'b000100110000111000001110;
rgb[34] = 24'b001001100001110100011101;
rgb[35] = 24'b001110010010110000101100;
rgb[36] = 24'b010011010011101000111010;
rgb[37] = 24'b011000000100100101001001;
rgb[38] = 24'b011100110101100001011000;
rgb[39] = 24'b100001100110011101100111;
rgb[40] = 24'b100101110111100001111000;
rgb[41] = 24'b101001101000101110001011;
rgb[42] = 24'b101101011001111010011110;
rgb[43] = 24'b110001001011000110110001;
rgb[44] = 24'b110100101100010111000101;
rgb[45] = 24'b111000011101100011011000;
rgb[46] = 24'b111100001110101111101011;
rgb[47] = 24'b111111111111111111111111;
rgb[48] = 24'b000000000000000000000000;
rgb[49] = 24'b000101000000110100001101;
rgb[50] = 24'b001010000001101100011011;
rgb[51] = 24'b001111010010100000101000;
rgb[52] = 24'b010100010011011000110110;
rgb[53] = 24'b011001010100010001000100;
rgb[54] = 24'b011110100101000101010001;
rgb[55] = 24'b100011100101111101011111;
rgb[56] = 24'b100111110111000001110000;
rgb[57] = 24'b101011011000010010000100;
rgb[58] = 24'b101110111001100010011000;
rgb[59] = 24'b110010001010110110101101;
rgb[60] = 24'b110101101100000111000001;
rgb[61] = 24'b111000111101011011010110;
rgb[62] = 24'b111100011110101011101010;
rgb[63] = 24'b111111111111111111111111;
rgb[64] = 24'b000000000000000000000000;
rgb[65] = 24'b000101010000110000001100;
rgb[66] = 24'b001010110001100000011000;
rgb[67] = 24'b010000000010010100100101;
rgb[68] = 24'b010101100011000100110001;
rgb[69] = 24'b011010110011111000111110;
rgb[70] = 24'b100000010100101001001010;
rgb[71] = 24'b100101100101011101010111;
rgb[72] = 24'b101001110110100001101000;
rgb[73] = 24'b101101000111110101111101;
rgb[74] = 24'b110000001001001110010011;
rgb[75] = 24'b110011011010100010101000;
rgb[76] = 24'b110110011011111010111110;
rgb[77] = 24'b111001101101001111010011;
rgb[78] = 24'b111100101110100111101001;
rgb[79] = 24'b111111111111111111111111;
rgb[80] = 24'b000000000000000000000000;
rgb[81] = 24'b000101100000101100001011;
rgb[82] = 24'b001011010001011000010110;
rgb[83] = 24'b010001000010001000100010;
rgb[84] = 24'b010110100010110100101101;
rgb[85] = 24'b011100010011100000111000;
rgb[86] = 24'b100010000100010001000100;
rgb[87] = 24'b100111100100111101001111;
rgb[88] = 24'b101011110110000001100000;
rgb[89] = 24'b101110110111011001110110;
rgb[90] = 24'b110001101000110110001101;
rgb[91] = 24'b110100011010010010100100;
rgb[92] = 24'b110111011011101110111011;
rgb[93] = 24'b111010001101000111010001;
rgb[94] = 24'b111100111110100011101000;
rgb[95] = 24'b111111111111111111111111;
rgb[96] = 24'b000000000000000000000000;
rgb[97] = 24'b000101110000101000001010;
rgb[98] = 24'b001011110001010000010100;
rgb[99] = 24'b010001110001111000011110;
rgb[100] = 24'b010111110010100000101000;
rgb[101] = 24'b011101100011001100110011;
rgb[102] = 24'b100011100011110100111101;
rgb[103] = 24'b101001100100011101000111;
rgb[104] = 24'b101101110101100001011000;
rgb[105] = 24'b110000010111000001110000;
rgb[106] = 24'b110011001000011110000111;
rgb[107] = 24'b110101101001111110011111;
rgb[108] = 24'b111000001011011110110111;
rgb[109] = 24'b111010101100111111001111;
rgb[110] = 24'b111101001110011111100111;
rgb[111] = 24'b111111101111111111111111;
rgb[112] = 24'b000000000000000000000000;
rgb[113] = 24'b000110000000100100001001;
rgb[114] = 24'b001100010001001000010010;
rgb[115] = 24'b010010100001101100011011;
rgb[116] = 24'b011000110010010000100100;
rgb[117] = 24'b011111000010110100101101;
rgb[118] = 24'b100101010011011000110110;
rgb[119] = 24'b101011100011111100111111;
rgb[120] = 24'b101111110101000001010000;
rgb[121] = 24'b110010000110100101101001;
rgb[122] = 24'b110100011000001010000010;
rgb[123] = 24'b110110101001101110011011;
rgb[124] = 24'b111000111011010010110100;
rgb[125] = 24'b111011001100110111001101;
rgb[126] = 24'b111101011110011011100110;
rgb[127] = 24'b111111111111111111111111;
rgb[128] = 24'b000000000000000000000000;
rgb[129] = 24'b000110100000011100000111;
rgb[130] = 24'b001101000000111100001111;
rgb[131] = 24'b010011100001011100010111;
rgb[132] = 24'b011010000001111100011111;
rgb[133] = 24'b100000100010011100100111;
rgb[134] = 24'b100111000010111100101111;
rgb[135] = 24'b101101100011011100110111;
rgb[136] = 24'b110001110100100001001000;
rgb[137] = 24'b110011110110001001100010;
rgb[138] = 24'b110101110111110001111100;
rgb[139] = 24'b110111111001011010010110;
rgb[140] = 24'b111001111011000010110000;
rgb[141] = 24'b111011111100101011001010;
rgb[142] = 24'b111101111110010011100100;
rgb[143] = 24'b111111101111111111111111;
rgb[144] = 24'b000000000000000000000000;
rgb[145] = 24'b000110110000011000000110;
rgb[146] = 24'b001101100000110100001101;
rgb[147] = 24'b010100010001010000010100;
rgb[148] = 24'b011011000001101100011011;
rgb[149] = 24'b100010000010000100100001;
rgb[150] = 24'b101000110010100000101000;
rgb[151] = 24'b101111100010111100101111;
rgb[152] = 24'b110011110100000001000000;
rgb[153] = 24'b110101100101101101011011;
rgb[154] = 24'b110111010111011001110110;
rgb[155] = 24'b111000111001001010010010;
rgb[156] = 24'b111010101010110110101101;
rgb[157] = 24'b111100011100100011001000;
rgb[158] = 24'b111110001110001111100011;
rgb[159] = 24'b111111111111111111111111;
rgb[160] = 24'b000000000000000000000000;
rgb[161] = 24'b000111000000010100000101;
rgb[162] = 24'b001110000000101100001011;
rgb[163] = 24'b010101010001000100010001;
rgb[164] = 24'b011100010001011000010110;
rgb[165] = 24'b100011010001110000011100;
rgb[166] = 24'b101010100010001000100010;
rgb[167] = 24'b110001100010011100100111;
rgb[168] = 24'b110101110011100000111000;
rgb[169] = 24'b110111010101010001010100;
rgb[170] = 24'b111000100111000101110001;
rgb[171] = 24'b111010001000110110001101;
rgb[172] = 24'b111011101010101010101010;
rgb[173] = 24'b111100111100011011000110;
rgb[174] = 24'b111110011110001011100010;
rgb[175] = 24'b111111101111111111111111;
rgb[176] = 24'b000000000000000000000000;
rgb[177] = 24'b000111010000010000000100;
rgb[178] = 24'b001110100000100100001001;
rgb[179] = 24'b010110000000110100001101;
rgb[180] = 24'b011101010001001000010010;
rgb[181] = 24'b100100110001011000010110;
rgb[182] = 24'b101100000001101100011011;
rgb[183] = 24'b110011100001111100011111;
rgb[184] = 24'b110111110011000000110000;
rgb[185] = 24'b111000110100111001001110;
rgb[186] = 24'b111010000110101101101011;
rgb[187] = 24'b111011001000100110001001;
rgb[188] = 24'b111100011010011010100110;
rgb[189] = 24'b111101011100010011000100;
rgb[190] = 24'b111110101110000111100001;
rgb[191] = 24'b111111111111111111111111;
rgb[192] = 24'b000000000000000000000000;
rgb[193] = 24'b000111100000001100000011;
rgb[194] = 24'b001111010000011000000110;
rgb[195] = 24'b010110110000101000001010;
rgb[196] = 24'b011110100000110100001101;
rgb[197] = 24'b100110010001000000010000;
rgb[198] = 24'b101101110001010000010100;
rgb[199] = 24'b110101100001011100010111;
rgb[200] = 24'b111001110010100000101000;
rgb[201] = 24'b111010100100011101000111;
rgb[202] = 24'b111011100110010101100101;
rgb[203] = 24'b111100011000010010000100;
rgb[204] = 24'b111101001010001110100011;
rgb[205] = 24'b111110001100000111000001;
rgb[206] = 24'b111110111110000011100000;
rgb[207] = 24'b111111111111111111111111;
rgb[208] = 24'b000000000000000000000000;
rgb[209] = 24'b000111110000001000000010;
rgb[210] = 24'b001111110000010000000100;
rgb[211] = 24'b010111110000011000000110;
rgb[212] = 24'b011111100000100100001001;
rgb[213] = 24'b100111100000101100001011;
rgb[214] = 24'b101111100000110100001101;
rgb[215] = 24'b110111100000111100001111;
rgb[216] = 24'b111011110010000000100000;
rgb[217] = 24'b111100010100000001000000;
rgb[218] = 24'b111100110110000001100000;
rgb[219] = 24'b111101011000000010000000;
rgb[220] = 24'b111110001001111110011111;
rgb[221] = 24'b111110101011111110111111;
rgb[222] = 24'b111111001101111111011111;
rgb[223] = 24'b111111111111111111111111;
rgb[224] = 24'b000000000000000000000000;
rgb[225] = 24'b001000000000000100000001;
rgb[226] = 24'b010000010000001000000010;
rgb[227] = 24'b011000100000001100000011;
rgb[228] = 24'b100000110000010000000100;
rgb[229] = 24'b101001000000010100000101;
rgb[230] = 24'b110001010000011000000110;
rgb[231] = 24'b111001100000011100000111;
rgb[232] = 24'b111101110001100000011000;
rgb[233] = 24'b111110000011100100111001;
rgb[234] = 24'b111110010101101001011010;
rgb[235] = 24'b111110100111101101111011;
rgb[236] = 24'b111110111001110010011100;
rgb[237] = 24'b111111001011110110111101;
rgb[238] = 24'b111111011101111011011110;
rgb[239] = 24'b111111111111111111111111;
rgb[240] = 24'b000000000000000000000000;
rgb[241] = 24'b001000100000000000000000;
rgb[242] = 24'b010001000000000000000000;
rgb[243] = 24'b011001100000000000000000;
rgb[244] = 24'b100010000000000000000000;
rgb[245] = 24'b101010100000000000000000;
rgb[246] = 24'b110011000000000000000000;
rgb[247] = 24'b111011100000000000000000;
rgb[248] = 24'b111111100001000100010001;
rgb[249] = 24'b111111110011001000110010;
rgb[250] = 24'b111111100101010101010101;
rgb[251] = 24'b111111110111011001110110;
rgb[252] = 24'b111111111001100110011001;
rgb[253] = 24'b111111111011101110111011;
rgb[254] = 24'b111111111101110111011101;
rgb[255] = 24'b111111111111111111111111;
rgb[256] = 24'b000000000000000000000000;
rgb[257] = 24'b000100010001000100010001;
rgb[258] = 24'b001000100010001000100010;
rgb[259] = 24'b001100110011001100110011;
rgb[260] = 24'b010001000100010001000100;
rgb[261] = 24'b010101010101010101010101;
rgb[262] = 24'b011001100110011001100110;
rgb[263] = 24'b011101110111011101110111;
rgb[264] = 24'b100010001000100010001000;
rgb[265] = 24'b100110011001100110011001;
rgb[266] = 24'b101010101010101010101010;
rgb[267] = 24'b101110111011101110111011;
rgb[268] = 24'b110011001100110011001100;
rgb[269] = 24'b110111011101110111011101;
rgb[270] = 24'b111011101110111011101110;
rgb[271] = 24'b111111111111111111111111;
rgb[272] = 24'b000000000000000000000000;
rgb[273] = 24'b000100100001000000001111;
rgb[274] = 24'b001001000010000000011111;
rgb[275] = 24'b001101100011000000101111;
rgb[276] = 24'b010010000100000000111111;
rgb[277] = 24'b010110100101000001001111;
rgb[278] = 24'b011011000110000001011111;
rgb[279] = 24'b011111100111000001101111;
rgb[280] = 24'b100011111000000110000000;
rgb[281] = 24'b100111111001001110010010;
rgb[282] = 24'b101011111010010110100100;
rgb[283] = 24'b101111111011011110110110;
rgb[284] = 24'b110011111100100111001000;
rgb[285] = 24'b110111111101101111011010;
rgb[286] = 24'b111011111110110111101100;
rgb[287] = 24'b111111111111111111111111;
rgb[288] = 24'b000000000000000000000000;
rgb[289] = 24'b000100110000111100001110;
rgb[290] = 24'b001001100001111000011101;
rgb[291] = 24'b001110010010110100101100;
rgb[292] = 24'b010011010011110000111010;
rgb[293] = 24'b011000000100101101001001;
rgb[294] = 24'b011100110101101001011000;
rgb[295] = 24'b100001100110101001100111;
rgb[296] = 24'b100101110111101101111000;
rgb[297] = 24'b101001101000110110001011;
rgb[298] = 24'b101101011010000010011110;
rgb[299] = 24'b110001001011001110110001;
rgb[300] = 24'b110100101100011011000101;
rgb[301] = 24'b111000011101100111011000;
rgb[302] = 24'b111100001110110011101011;
rgb[303] = 24'b111111111111111111111111;
rgb[304] = 24'b000000000000000000000000;
rgb[305] = 24'b000101000000111000001101;
rgb[306] = 24'b001010000001110000011011;
rgb[307] = 24'b001111010010101000101000;
rgb[308] = 24'b010100010011100000110110;
rgb[309] = 24'b011001010100011101000100;
rgb[310] = 24'b011110100101010101010001;
rgb[311] = 24'b100011100110001101011111;
rgb[312] = 24'b100111110111010001110000;
rgb[313] = 24'b101011011000100010000100;
rgb[314] = 24'b101110111001110010011000;
rgb[315] = 24'b110010001010111110101101;
rgb[316] = 24'b110101101100001111000001;
rgb[317] = 24'b111000111101011111010110;
rgb[318] = 24'b111100011110101111101010;
rgb[319] = 24'b111111111111111111111111;
rgb[320] = 24'b000000000000000000000000;
rgb[321] = 24'b000101010000110100001100;
rgb[322] = 24'b001010110001101000011000;
rgb[323] = 24'b010000000010011100100101;
rgb[324] = 24'b010101100011010100110001;
rgb[325] = 24'b011010110100001000111110;
rgb[326] = 24'b100000010100111101001010;
rgb[327] = 24'b100101100101110101010111;
rgb[328] = 24'b101001110110111001101000;
rgb[329] = 24'b101101001000001001111101;
rgb[330] = 24'b110000001001011110010011;
rgb[331] = 24'b110011011010110010101000;
rgb[332] = 24'b110110011100000010111110;
rgb[333] = 24'b111001101101010111010011;
rgb[334] = 24'b111100101110101011101001;
rgb[335] = 24'b111111111111111111111111;
rgb[336] = 24'b000000000000000000000000;
rgb[337] = 24'b000101100000110000001011;
rgb[338] = 24'b001011010001100000010110;
rgb[339] = 24'b010001000010010100100010;
rgb[340] = 24'b010110100011000100101101;
rgb[341] = 24'b011100010011111000111000;
rgb[342] = 24'b100010000100101001000100;
rgb[343] = 24'b100111100101011001001111;
rgb[344] = 24'b101011110110011101100000;
rgb[345] = 24'b101110110111110101110110;
rgb[346] = 24'b110001101001001110001101;
rgb[347] = 24'b110100011010100010100100;
rgb[348] = 24'b110111011011111010111011;
rgb[349] = 24'b111010001101001111010001;
rgb[350] = 24'b111100111110100111101000;
rgb[351] = 24'b111111111111111111111111;
rgb[352] = 24'b000000000000000000000000;
rgb[353] = 24'b000101110000101100001010;
rgb[354] = 24'b001011110001011000010100;
rgb[355] = 24'b010001110010001000011110;
rgb[356] = 24'b010111110010110100101000;
rgb[357] = 24'b011101100011100100110011;
rgb[358] = 24'b100011100100010000111101;
rgb[359] = 24'b101001100101000001000111;
rgb[360] = 24'b101101110110000101011000;
rgb[361] = 24'b110000010111011101110000;
rgb[362] = 24'b110011001000111010000111;
rgb[363] = 24'b110101101010010010011111;
rgb[364] = 24'b111000001011101110110111;
rgb[365] = 24'b111010101101000111001111;
rgb[366] = 24'b111101001110100011100111;
rgb[367] = 24'b111111101111111111111111;
rgb[368] = 24'b000000000000000000000000;
rgb[369] = 24'b000110000000101000001001;
rgb[370] = 24'b001100010001010100010010;
rgb[371] = 24'b010010100001111100011011;
rgb[372] = 24'b011000110010101000100100;
rgb[373] = 24'b011111000011010000101101;
rgb[374] = 24'b100101010011111100110110;
rgb[375] = 24'b101011100100101000111111;
rgb[376] = 24'b101111110101101101010000;
rgb[377] = 24'b110010000111001001101001;
rgb[378] = 24'b110100011000100110000010;
rgb[379] = 24'b110110101010000110011011;
rgb[380] = 24'b111000111011100010110100;
rgb[381] = 24'b111011001101000011001101;
rgb[382] = 24'b111101011110011111100110;
rgb[383] = 24'b111111111111111111111111;
rgb[384] = 24'b000000000000000000000000;
rgb[385] = 24'b000110100000100100000111;
rgb[386] = 24'b001101000001001100001111;
rgb[387] = 24'b010011100001110000010111;
rgb[388] = 24'b011010000010011000011111;
rgb[389] = 24'b100000100011000000100111;
rgb[390] = 24'b100111000011100100101111;
rgb[391] = 24'b101101100100001100110111;
rgb[392] = 24'b110001110101010001001000;
rgb[393] = 24'b110011110110110001100010;
rgb[394] = 24'b110101111000010101111100;
rgb[395] = 24'b110111111001110110010110;
rgb[396] = 24'b111001111011010110110000;
rgb[397] = 24'b111011111100111011001010;
rgb[398] = 24'b111101111110011011100100;
rgb[399] = 24'b111111101111111111111111;
rgb[400] = 24'b000000000000000000000000;
rgb[401] = 24'b000110110000100000000110;
rgb[402] = 24'b001101100001000100001101;
rgb[403] = 24'b010100010001101000010100;
rgb[404] = 24'b011011000010001000011011;
rgb[405] = 24'b100010000010101100100001;
rgb[406] = 24'b101000110011010000101000;
rgb[407] = 24'b101111100011110100101111;
rgb[408] = 24'b110011110100111001000000;
rgb[409] = 24'b110101100110011101011011;
rgb[410] = 24'b110111011000000001110110;
rgb[411] = 24'b111000111001100110010010;
rgb[412] = 24'b111010101011001110101101;
rgb[413] = 24'b111100011100110011001000;
rgb[414] = 24'b111110001110010111100011;
rgb[415] = 24'b111111111111111111111111;
rgb[416] = 24'b000000000000000000000000;
rgb[417] = 24'b000111000000011100000101;
rgb[418] = 24'b001110000000111100001011;
rgb[419] = 24'b010101010001011100010001;
rgb[420] = 24'b011100010001111100010110;
rgb[421] = 24'b100011010010011100011100;
rgb[422] = 24'b101010100010111000100010;
rgb[423] = 24'b110001100011011000100111;
rgb[424] = 24'b110101110100011100111000;
rgb[425] = 24'b110111010110000101010100;
rgb[426] = 24'b111000100111110001110001;
rgb[427] = 24'b111010001001011010001101;
rgb[428] = 24'b111011101011000010101010;
rgb[429] = 24'b111100111100101011000110;
rgb[430] = 24'b111110011110010011100010;
rgb[431] = 24'b111111101111111111111111;
rgb[432] = 24'b000000000000000000000000;
rgb[433] = 24'b000111010000011000000100;
rgb[434] = 24'b001110100000110100001001;
rgb[435] = 24'b010110000001010000001101;
rgb[436] = 24'b011101010001101100010010;
rgb[437] = 24'b100100110010001000010110;
rgb[438] = 24'b101100000010100100011011;
rgb[439] = 24'b110011100011000000011111;
rgb[440] = 24'b110111110100000100110000;
rgb[441] = 24'b111000110101110001001110;
rgb[442] = 24'b111010000111011101101011;
rgb[443] = 24'b111011001001001010001001;
rgb[444] = 24'b111100011010110110100110;
rgb[445] = 24'b111101011100100011000100;
rgb[446] = 24'b111110101110001111100001;
rgb[447] = 24'b111111111111111111111111;
rgb[448] = 24'b000000000000000000000000;
rgb[449] = 24'b000111100000010100000011;
rgb[450] = 24'b001111010000101100000110;
rgb[451] = 24'b010110110001000100001010;
rgb[452] = 24'b011110100001011100001101;
rgb[453] = 24'b100110010001110100010000;
rgb[454] = 24'b101101110010001100010100;
rgb[455] = 24'b110101100010100100010111;
rgb[456] = 24'b111001110011101000101000;
rgb[457] = 24'b111010100101011001000111;
rgb[458] = 24'b111011100111001001100101;
rgb[459] = 24'b111100011000111010000100;
rgb[460] = 24'b111101001010101010100011;
rgb[461] = 24'b111110001100011011000001;
rgb[462] = 24'b111110111110001011100000;
rgb[463] = 24'b111111111111111111111111;
rgb[464] = 24'b000000000000000000000000;
rgb[465] = 24'b000111110000010100000010;
rgb[466] = 24'b001111110000101000000100;
rgb[467] = 24'b010111110000111100000110;
rgb[468] = 24'b011111100001010000001001;
rgb[469] = 24'b100111100001100100001011;
rgb[470] = 24'b101111100001111000001101;
rgb[471] = 24'b110111100010001100001111;
rgb[472] = 24'b111011110011010000100000;
rgb[473] = 24'b111100010101000101000000;
rgb[474] = 24'b111100110110111001100000;
rgb[475] = 24'b111101011000101110000000;
rgb[476] = 24'b111110001010100010011111;
rgb[477] = 24'b111110101100010110111111;
rgb[478] = 24'b111111001110001011011111;
rgb[479] = 24'b111111111111111111111111;
rgb[480] = 24'b000000000000000000000000;
rgb[481] = 24'b001000000000010000000001;
rgb[482] = 24'b010000010000100000000010;
rgb[483] = 24'b011000100000110000000011;
rgb[484] = 24'b100000110001000000000100;
rgb[485] = 24'b101001000001010000000101;
rgb[486] = 24'b110001010001100000000110;
rgb[487] = 24'b111001100001110100000111;
rgb[488] = 24'b111101110010111000011000;
rgb[489] = 24'b111110000100101100111001;
rgb[490] = 24'b111110010110100101011010;
rgb[491] = 24'b111110101000011101111011;
rgb[492] = 24'b111110111010010110011100;
rgb[493] = 24'b111111001100001110111101;
rgb[494] = 24'b111111011110000111011110;
rgb[495] = 24'b111111111111111111111111;
rgb[496] = 24'b000000000000000000000000;
rgb[497] = 24'b001000100000001100000000;
rgb[498] = 24'b010001000000011000000000;
rgb[499] = 24'b011001100000100100000000;
rgb[500] = 24'b100010000000110000000000;
rgb[501] = 24'b101010100001000000000000;
rgb[502] = 24'b110011000001001100000000;
rgb[503] = 24'b111011100001011000000000;
rgb[504] = 24'b111111100010011100010001;
rgb[505] = 24'b111111110100011000110010;
rgb[506] = 24'b111111100110010101010101;
rgb[507] = 24'b111111111000001101110110;
rgb[508] = 24'b111111111010001010011001;
rgb[509] = 24'b111111111100000110111011;
rgb[510] = 24'b111111111110000011011101;
rgb[511] = 24'b111111111111111111111111;
rgb[512] = 24'b000000000000000000000000;
rgb[513] = 24'b000100010001000100010001;
rgb[514] = 24'b001000100010001000100010;
rgb[515] = 24'b001100110011001100110011;
rgb[516] = 24'b010001000100010001000100;
rgb[517] = 24'b010101010101010101010101;
rgb[518] = 24'b011001100110011001100110;
rgb[519] = 24'b011101110111011101110111;
rgb[520] = 24'b100010001000100010001000;
rgb[521] = 24'b100110011001100110011001;
rgb[522] = 24'b101010101010101010101010;
rgb[523] = 24'b101110111011101110111011;
rgb[524] = 24'b110011001100110011001100;
rgb[525] = 24'b110111011101110111011101;
rgb[526] = 24'b111011101110111011101110;
rgb[527] = 24'b111111111111111111111111;
rgb[528] = 24'b000000000000000000000000;
rgb[529] = 24'b000100100001000000001111;
rgb[530] = 24'b001001000010000000011111;
rgb[531] = 24'b001101100011000000101111;
rgb[532] = 24'b010010000100000100111111;
rgb[533] = 24'b010110100101000101001111;
rgb[534] = 24'b011011000110000101011111;
rgb[535] = 24'b011111100111001001101111;
rgb[536] = 24'b100011111000001110000000;
rgb[537] = 24'b100111111001010010010010;
rgb[538] = 24'b101011111010011010100100;
rgb[539] = 24'b101111111011100010110110;
rgb[540] = 24'b110011111100100111001000;
rgb[541] = 24'b110111111101101111011010;
rgb[542] = 24'b111011111110110111101100;
rgb[543] = 24'b111111111111111111111111;
rgb[544] = 24'b000000000000000000000000;
rgb[545] = 24'b000100110000111100001110;
rgb[546] = 24'b001001100001111100011101;
rgb[547] = 24'b001110010010111000101100;
rgb[548] = 24'b010011010011111000111010;
rgb[549] = 24'b011000000100110101001001;
rgb[550] = 24'b011100110101110101011000;
rgb[551] = 24'b100001100110110101100111;
rgb[552] = 24'b100101110111111001111000;
rgb[553] = 24'b101001101001000010001011;
rgb[554] = 24'b101101011010001010011110;
rgb[555] = 24'b110001001011010110110001;
rgb[556] = 24'b110100101100011111000101;
rgb[557] = 24'b111000011101101011011000;
rgb[558] = 24'b111100001110110011101011;
rgb[559] = 24'b111111111111111111111111;
rgb[560] = 24'b000000000000000000000000;
rgb[561] = 24'b000101000000111000001101;
rgb[562] = 24'b001010000001110100011011;
rgb[563] = 24'b001111010010110000101000;
rgb[564] = 24'b010100010011101100110110;
rgb[565] = 24'b011001010100101001000100;
rgb[566] = 24'b011110100101100101010001;
rgb[567] = 24'b100011100110100001011111;
rgb[568] = 24'b100111110111100101110000;
rgb[569] = 24'b101011011000110010000100;
rgb[570] = 24'b101110111001111110011000;
rgb[571] = 24'b110010001011001010101101;
rgb[572] = 24'b110101101100010111000001;
rgb[573] = 24'b111000111101100011010110;
rgb[574] = 24'b111100011110101111101010;
rgb[575] = 24'b111111111111111111111111;
rgb[576] = 24'b000000000000000000000000;
rgb[577] = 24'b000101010000111000001100;
rgb[578] = 24'b001010110001110000011000;
rgb[579] = 24'b010000000010101000100101;
rgb[580] = 24'b010101100011100000110001;
rgb[581] = 24'b011010110100011000111110;
rgb[582] = 24'b100000010101010101001010;
rgb[583] = 24'b100101100110001101010111;
rgb[584] = 24'b101001110111010001101000;
rgb[585] = 24'b101101001000100001111101;
rgb[586] = 24'b110000001001101110010011;
rgb[587] = 24'b110011011010111110101000;
rgb[588] = 24'b110110011100001110111110;
rgb[589] = 24'b111001101101011111010011;
rgb[590] = 24'b111100101110101111101001;
rgb[591] = 24'b111111111111111111111111;
rgb[592] = 24'b000000000000000000000000;
rgb[593] = 24'b000101100000110100001011;
rgb[594] = 24'b001011010001101000010110;
rgb[595] = 24'b010001000010100000100010;
rgb[596] = 24'b010110100011010100101101;
rgb[597] = 24'b011100010100001100111000;
rgb[598] = 24'b100010000101000001000100;
rgb[599] = 24'b100111100101111001001111;
rgb[600] = 24'b101011110110111101100000;
rgb[601] = 24'b101110111000001101110110;
rgb[602] = 24'b110001101001100010001101;
rgb[603] = 24'b110100011010110010100100;
rgb[604] = 24'b110111011100000110111011;
rgb[605] = 24'b111010001101010111010001;
rgb[606] = 24'b111100111110101011101000;
rgb[607] = 24'b111111111111111111111111;
rgb[608] = 24'b000000000000000000000000;
rgb[609] = 24'b000101110000110000001010;
rgb[610] = 24'b001011110001100100010100;
rgb[611] = 24'b010001110010011000011110;
rgb[612] = 24'b010111110011001100101000;
rgb[613] = 24'b011101100011111100110011;
rgb[614] = 24'b100011100100110000111101;
rgb[615] = 24'b101001100101100101000111;
rgb[616] = 24'b101101110110101001011000;
rgb[617] = 24'b110000010111111101110000;
rgb[618] = 24'b110011001001010010000111;
rgb[619] = 24'b110101101010101010011111;
rgb[620] = 24'b111000001011111110110111;
rgb[621] = 24'b111010101101010011001111;
rgb[622] = 24'b111101001110100111100111;
rgb[623] = 24'b111111101111111111111111;
rgb[624] = 24'b000000000000000000000000;
rgb[625] = 24'b000110000000110000001001;
rgb[626] = 24'b001100010001100000010010;
rgb[627] = 24'b010010100010010000011011;
rgb[628] = 24'b011000110011000000100100;
rgb[629] = 24'b011111000011110000101101;
rgb[630] = 24'b100101010100100000110110;
rgb[631] = 24'b101011100101010000111111;
rgb[632] = 24'b101111110110010101010000;
rgb[633] = 24'b110010000111101101101001;
rgb[634] = 24'b110100011001000110000010;
rgb[635] = 24'b110110101010011110011011;
rgb[636] = 24'b111000111011110110110100;
rgb[637] = 24'b111011001101001111001101;
rgb[638] = 24'b111101011110100111100110;
rgb[639] = 24'b111111111111111111111111;
rgb[640] = 24'b000000000000000000000000;
rgb[641] = 24'b000110100000101100000111;
rgb[642] = 24'b001101000001011000001111;
rgb[643] = 24'b010011100010001000010111;
rgb[644] = 24'b011010000010110100011111;
rgb[645] = 24'b100000100011100000100111;
rgb[646] = 24'b100111000100010000101111;
rgb[647] = 24'b101101100100111100110111;
rgb[648] = 24'b110001110110000001001000;
rgb[649] = 24'b110011110111011101100010;
rgb[650] = 24'b110101111000110101111100;
rgb[651] = 24'b110111111010010010010110;
rgb[652] = 24'b111001111011101110110000;
rgb[653] = 24'b111011111101000111001010;
rgb[654] = 24'b111101111110100011100100;
rgb[655] = 24'b111111101111111111111111;
rgb[656] = 24'b000000000000000000000000;
rgb[657] = 24'b000110110000101000000110;
rgb[658] = 24'b001101100001010100001101;
rgb[659] = 24'b010100010010000000010100;
rgb[660] = 24'b011011000010101000011011;
rgb[661] = 24'b100010000011010100100001;
rgb[662] = 24'b101000110100000000101000;
rgb[663] = 24'b101111100100101000101111;
rgb[664] = 24'b110011110101101101000000;
rgb[665] = 24'b110101100111001101011011;
rgb[666] = 24'b110111011000101001110110;
rgb[667] = 24'b111000111010000110010010;
rgb[668] = 24'b111010101011100110101101;
rgb[669] = 24'b111100011101000011001000;
rgb[670] = 24'b111110001110011111100011;
rgb[671] = 24'b111111111111111111111111;
rgb[672] = 24'b000000000000000000000000;
rgb[673] = 24'b000111000000100100000101;
rgb[674] = 24'b001110000001001100001011;
rgb[675] = 24'b010101010001110100010001;
rgb[676] = 24'b011100010010011100010110;
rgb[677] = 24'b100011010011000100011100;
rgb[678] = 24'b101010100011101100100010;
rgb[679] = 24'b110001100100010100100111;
rgb[680] = 24'b110101110101011000111000;
rgb[681] = 24'b110111010110111001010100;
rgb[682] = 24'b111000101000011001110001;
rgb[683] = 24'b111010001001111010001101;
rgb[684] = 24'b111011101011011010101010;
rgb[685] = 24'b111100111100111011000110;
rgb[686] = 24'b111110011110011011100010;
rgb[687] = 24'b111111101111111111111111;
rgb[688] = 24'b000000000000000000000000;
rgb[689] = 24'b000111010000100100000100;
rgb[690] = 24'b001110100001001000001001;
rgb[691] = 24'b010110000001101100001101;
rgb[692] = 24'b011101010010010100010010;
rgb[693] = 24'b100100110010111000010110;
rgb[694] = 24'b101100000011011100011011;
rgb[695] = 24'b110011100100000000011111;
rgb[696] = 24'b110111110101000100110000;
rgb[697] = 24'b111000110110101001001110;
rgb[698] = 24'b111010001000001101101011;
rgb[699] = 24'b111011001001110010001001;
rgb[700] = 24'b111100011011010010100110;
rgb[701] = 24'b111101011100110111000100;
rgb[702] = 24'b111110101110011011100001;
rgb[703] = 24'b111111111111111111111111;
rgb[704] = 24'b000000000000000000000000;
rgb[705] = 24'b000111100000100000000011;
rgb[706] = 24'b001111010001000100000110;
rgb[707] = 24'b010110110001100100001010;
rgb[708] = 24'b011110100010001000001101;
rgb[709] = 24'b100110010010101000010000;
rgb[710] = 24'b101101110011001100010100;
rgb[711] = 24'b110101100011110000010111;
rgb[712] = 24'b111001110100110100101000;
rgb[713] = 24'b111010100110011001000111;
rgb[714] = 24'b111011100111111101100101;
rgb[715] = 24'b111100011001100110000100;
rgb[716] = 24'b111101001011001010100011;
rgb[717] = 24'b111110001100110011000001;
rgb[718] = 24'b111110111110010111100000;
rgb[719] = 24'b111111111111111111111111;
rgb[720] = 24'b000000000000000000000000;
rgb[721] = 24'b000111110000011100000010;
rgb[722] = 24'b001111110000111100000100;
rgb[723] = 24'b010111110001011100000110;
rgb[724] = 24'b011111100001111100001001;
rgb[725] = 24'b100111100010011100001011;
rgb[726] = 24'b101111100010111100001101;
rgb[727] = 24'b110111100011011100001111;
rgb[728] = 24'b111011110100100000100000;
rgb[729] = 24'b111100010110001001000000;
rgb[730] = 24'b111100110111110001100000;
rgb[731] = 24'b111101011001011010000000;
rgb[732] = 24'b111110001011000010011111;
rgb[733] = 24'b111110101100101010111111;
rgb[734] = 24'b111111001110010011011111;
rgb[735] = 24'b111111111111111111111111;
rgb[736] = 24'b000000000000000000000000;
rgb[737] = 24'b001000000000011100000001;
rgb[738] = 24'b010000010000111000000010;
rgb[739] = 24'b011000100001010100000011;
rgb[740] = 24'b100000110001110000000100;
rgb[741] = 24'b101001000010001100000101;
rgb[742] = 24'b110001010010101100000110;
rgb[743] = 24'b111001100011001000000111;
rgb[744] = 24'b111101110100001100011000;
rgb[745] = 24'b111110000101111000111001;
rgb[746] = 24'b111110010111100001011010;
rgb[747] = 24'b111110101001001101111011;
rgb[748] = 24'b111110111010111010011100;
rgb[749] = 24'b111111001100100110111101;
rgb[750] = 24'b111111011110010011011110;
rgb[751] = 24'b111111111111111111111111;
rgb[752] = 24'b000000000000000000000000;
rgb[753] = 24'b001000100000011000000000;
rgb[754] = 24'b010001000000110000000000;
rgb[755] = 24'b011001100001001100000000;
rgb[756] = 24'b100010000001100100000000;
rgb[757] = 24'b101010100010000000000000;
rgb[758] = 24'b110011000010011000000000;
rgb[759] = 24'b111011100010110100000000;
rgb[760] = 24'b111111100011111000010001;
rgb[761] = 24'b111111110101100100110010;
rgb[762] = 24'b111111100111010101010101;
rgb[763] = 24'b111111111001000001110110;
rgb[764] = 24'b111111111010110010011001;
rgb[765] = 24'b111111111100011110111011;
rgb[766] = 24'b111111111110001111011101;
rgb[767] = 24'b111111111111111111111111;
rgb[768] = 24'b000000000000000000000000;
rgb[769] = 24'b000100010001000100010001;
rgb[770] = 24'b001000100010001000100010;
rgb[771] = 24'b001100110011001100110011;
rgb[772] = 24'b010001000100010001000100;
rgb[773] = 24'b010101010101010101010101;
rgb[774] = 24'b011001100110011001100110;
rgb[775] = 24'b011101110111011101110111;
rgb[776] = 24'b100010001000100010001000;
rgb[777] = 24'b100110011001100110011001;
rgb[778] = 24'b101010101010101010101010;
rgb[779] = 24'b101110111011101110111011;
rgb[780] = 24'b110011001100110011001100;
rgb[781] = 24'b110111011101110111011101;
rgb[782] = 24'b111011101110111011101110;
rgb[783] = 24'b111111111111111111111111;
rgb[784] = 24'b000000000000000000000000;
rgb[785] = 24'b000100100001000000001111;
rgb[786] = 24'b001001000010000100011111;
rgb[787] = 24'b001101100011000100101111;
rgb[788] = 24'b010010000100001000111111;
rgb[789] = 24'b010110100101001001001111;
rgb[790] = 24'b011011000110001101011111;
rgb[791] = 24'b011111100111001101101111;
rgb[792] = 24'b100011111000010010000000;
rgb[793] = 24'b100111111001011010010010;
rgb[794] = 24'b101011111010011110100100;
rgb[795] = 24'b101111111011100110110110;
rgb[796] = 24'b110011111100101011001000;
rgb[797] = 24'b110111111101110011011010;
rgb[798] = 24'b111011111110110111101100;
rgb[799] = 24'b111111111111111111111111;
rgb[800] = 24'b000000000000000000000000;
rgb[801] = 24'b000100110001000000001110;
rgb[802] = 24'b001001100010000000011101;
rgb[803] = 24'b001110010011000000101100;
rgb[804] = 24'b010011010100000000111010;
rgb[805] = 24'b011000000101000001001001;
rgb[806] = 24'b011100110110000001011000;
rgb[807] = 24'b100001100111000001100111;
rgb[808] = 24'b100101111000000101111000;
rgb[809] = 24'b101001101001001110001011;
rgb[810] = 24'b101101011010010110011110;
rgb[811] = 24'b110001001011011110110001;
rgb[812] = 24'b110100101100100111000101;
rgb[813] = 24'b111000011101101111011000;
rgb[814] = 24'b111100001110110111101011;
rgb[815] = 24'b111111111111111111111111;
rgb[816] = 24'b000000000000000000000000;
rgb[817] = 24'b000101000000111100001101;
rgb[818] = 24'b001010000001111100011011;
rgb[819] = 24'b001111010010111000101000;
rgb[820] = 24'b010100010011111000110110;
rgb[821] = 24'b011001010100110101000100;
rgb[822] = 24'b011110100101110101010001;
rgb[823] = 24'b100011100110110001011111;
rgb[824] = 24'b100111110111110101110000;
rgb[825] = 24'b101011011001000010000100;
rgb[826] = 24'b101110111010001010011000;
rgb[827] = 24'b110010001011010110101101;
rgb[828] = 24'b110101101100011111000001;
rgb[829] = 24'b111000111101101011010110;
rgb[830] = 24'b111100011110110011101010;
rgb[831] = 24'b111111111111111111111111;
rgb[832] = 24'b000000000000000000000000;
rgb[833] = 24'b000101010000111100001100;
rgb[834] = 24'b001010110001111000011000;
rgb[835] = 24'b010000000010110100100101;
rgb[836] = 24'b010101100011110000110001;
rgb[837] = 24'b011010110100101100111110;
rgb[838] = 24'b100000010101101001001010;
rgb[839] = 24'b100101100110100101010111;
rgb[840] = 24'b101001110111101001101000;
rgb[841] = 24'b101101001000110101111101;
rgb[842] = 24'b110000001010000010010011;
rgb[843] = 24'b110011011011001110101000;
rgb[844] = 24'b110110011100011010111110;
rgb[845] = 24'b111001101101100111010011;
rgb[846] = 24'b111100101110110011101001;
rgb[847] = 24'b111111111111111111111111;
rgb[848] = 24'b000000000000000000000000;
rgb[849] = 24'b000101100000111000001011;
rgb[850] = 24'b001011010001110100010110;
rgb[851] = 24'b010001000010101100100010;
rgb[852] = 24'b010110100011101000101101;
rgb[853] = 24'b011100010100100000111000;
rgb[854] = 24'b100010000101011101000100;
rgb[855] = 24'b100111100110011001001111;
rgb[856] = 24'b101011110111011101100000;
rgb[857] = 24'b101110111000101001110110;
rgb[858] = 24'b110001101001110110001101;
rgb[859] = 24'b110100011011000110100100;
rgb[860] = 24'b110111011100010010111011;
rgb[861] = 24'b111010001101100011010001;
rgb[862] = 24'b111100111110101111101000;
rgb[863] = 24'b111111111111111111111111;
rgb[864] = 24'b000000000000000000000000;
rgb[865] = 24'b000101110000111000001010;
rgb[866] = 24'b001011110001110000010100;
rgb[867] = 24'b010001110010101000011110;
rgb[868] = 24'b010111110011100000101000;
rgb[869] = 24'b011101100100011000110011;
rgb[870] = 24'b100011100101010000111101;
rgb[871] = 24'b101001100110001001000111;
rgb[872] = 24'b101101110111001101011000;
rgb[873] = 24'b110000011000011101110000;
rgb[874] = 24'b110011001001101110000111;
rgb[875] = 24'b110101101010111110011111;
rgb[876] = 24'b111000001100001110110111;
rgb[877] = 24'b111010101101011111001111;
rgb[878] = 24'b111101001110101111100111;
rgb[879] = 24'b111111101111111111111111;
rgb[880] = 24'b000000000000000000000000;
rgb[881] = 24'b000110000000110100001001;
rgb[882] = 24'b001100010001101100010010;
rgb[883] = 24'b010010100010100000011011;
rgb[884] = 24'b011000110011011000100100;
rgb[885] = 24'b011111000100001100101101;
rgb[886] = 24'b100101010101000100110110;
rgb[887] = 24'b101011100101111100111111;
rgb[888] = 24'b101111110111000001010000;
rgb[889] = 24'b110010001000010001101001;
rgb[890] = 24'b110100011001100110000010;
rgb[891] = 24'b110110101010110110011011;
rgb[892] = 24'b111000111100000110110100;
rgb[893] = 24'b111011001101011011001101;
rgb[894] = 24'b111101011110101011100110;
rgb[895] = 24'b111111111111111111111111;
rgb[896] = 24'b000000000000000000000000;
rgb[897] = 24'b000110100000110100000111;
rgb[898] = 24'b001101000001101000001111;
rgb[899] = 24'b010011100010011100010111;
rgb[900] = 24'b011010000011010000011111;
rgb[901] = 24'b100000100100000100100111;
rgb[902] = 24'b100111000100111000101111;
rgb[903] = 24'b101101100101101100110111;
rgb[904] = 24'b110001110110110001001000;
rgb[905] = 24'b110011111000000101100010;
rgb[906] = 24'b110101111001011001111100;
rgb[907] = 24'b110111111010101110010110;
rgb[908] = 24'b111001111100000010110000;
rgb[909] = 24'b111011111101010111001010;
rgb[910] = 24'b111101111110101011100100;
rgb[911] = 24'b111111101111111111111111;
rgb[912] = 24'b000000000000000000000000;
rgb[913] = 24'b000110110000110000000110;
rgb[914] = 24'b001101100001100100001101;
rgb[915] = 24'b010100010010010100010100;
rgb[916] = 24'b011011000011001000011011;
rgb[917] = 24'b100010000011111100100001;
rgb[918] = 24'b101000110100101100101000;
rgb[919] = 24'b101111100101100000101111;
rgb[920] = 24'b110011110110100101000000;
rgb[921] = 24'b110101100111111001011011;
rgb[922] = 24'b110111011001010001110110;
rgb[923] = 24'b111000111010100110010010;
rgb[924] = 24'b111010101011111010101101;
rgb[925] = 24'b111100011101010011001000;
rgb[926] = 24'b111110001110100111100011;
rgb[927] = 24'b111111111111111111111111;
rgb[928] = 24'b000000000000000000000000;
rgb[929] = 24'b000111000000110000000101;
rgb[930] = 24'b001110000001100000001011;
rgb[931] = 24'b010101010010010000010001;
rgb[932] = 24'b011100010011000000010110;
rgb[933] = 24'b100011010011110000011100;
rgb[934] = 24'b101010100100100000100010;
rgb[935] = 24'b110001100101010100100111;
rgb[936] = 24'b110101110110010100111000;
rgb[937] = 24'b110111010111101101010100;
rgb[938] = 24'b111000101001000101110001;
rgb[939] = 24'b111010001010011110001101;
rgb[940] = 24'b111011101011110110101010;
rgb[941] = 24'b111100111101001111000110;
rgb[942] = 24'b111110011110100111100010;
rgb[943] = 24'b111111101111111111111111;
rgb[944] = 24'b000000000000000000000000;
rgb[945] = 24'b000111010000101100000100;
rgb[946] = 24'b001110100001011100001001;
rgb[947] = 24'b010110000010001000001101;
rgb[948] = 24'b011101010010111000010010;
rgb[949] = 24'b100100110011101000010110;
rgb[950] = 24'b101100000100010100011011;
rgb[951] = 24'b110011100101000100011111;
rgb[952] = 24'b110111110110001000110000;
rgb[953] = 24'b111000110111100001001110;
rgb[954] = 24'b111010001000111101101011;
rgb[955] = 24'b111011001010010110001001;
rgb[956] = 24'b111100011011101110100110;
rgb[957] = 24'b111101011101001011000100;
rgb[958] = 24'b111110101110100011100001;
rgb[959] = 24'b111111111111111111111111;
rgb[960] = 24'b000000000000000000000000;
rgb[961] = 24'b000111100000101100000011;
rgb[962] = 24'b001111010001011000000110;
rgb[963] = 24'b010110110010000100001010;
rgb[964] = 24'b011110100010110000001101;
rgb[965] = 24'b100110010011011100010000;
rgb[966] = 24'b101101110100001100010100;
rgb[967] = 24'b110101100100111000010111;
rgb[968] = 24'b111001110101111100101000;
rgb[969] = 24'b111010100111011001000111;
rgb[970] = 24'b111011101000110001100101;
rgb[971] = 24'b111100011010001110000100;
rgb[972] = 24'b111101001011101010100011;
rgb[973] = 24'b111110001101000111000001;
rgb[974] = 24'b111110111110100011100000;
rgb[975] = 24'b111111111111111111111111;
rgb[976] = 24'b000000000000000000000000;
rgb[977] = 24'b000111110000101000000010;
rgb[978] = 24'b001111110001010100000100;
rgb[979] = 24'b010111110010000000000110;
rgb[980] = 24'b011111100010101000001001;
rgb[981] = 24'b100111100011010100001011;
rgb[982] = 24'b101111100100000000001101;
rgb[983] = 24'b110111100100101000001111;
rgb[984] = 24'b111011110101101100100000;
rgb[985] = 24'b111100010111001101000000;
rgb[986] = 24'b111100111000101001100000;
rgb[987] = 24'b111101011010000110000000;
rgb[988] = 24'b111110001011100110011111;
rgb[989] = 24'b111110101101000010111111;
rgb[990] = 24'b111111001110011111011111;
rgb[991] = 24'b111111111111111111111111;
rgb[992] = 24'b000000000000000000000000;
rgb[993] = 24'b001000000000101000000001;
rgb[994] = 24'b010000010001010000000010;
rgb[995] = 24'b011000100001111000000011;
rgb[996] = 24'b100000110010100000000100;
rgb[997] = 24'b101001000011001100000101;
rgb[998] = 24'b110001010011110100000110;
rgb[999] = 24'b111001100100011100000111;
rgb[1000] = 24'b111101110101100000011000;
rgb[1001] = 24'b111110000111000000111001;
rgb[1002] = 24'b111110011000011101011010;
rgb[1003] = 24'b111110101001111101111011;
rgb[1004] = 24'b111110111011011110011100;
rgb[1005] = 24'b111111001100111110111101;
rgb[1006] = 24'b111111011110011111011110;
rgb[1007] = 24'b111111111111111111111111;
rgb[1008] = 24'b000000000000000000000000;
rgb[1009] = 24'b001000100000100100000000;
rgb[1010] = 24'b010001000001001100000000;
rgb[1011] = 24'b011001100001110100000000;
rgb[1012] = 24'b100010000010011000000000;
rgb[1013] = 24'b101010100011000000000000;
rgb[1014] = 24'b110011000011101000000000;
rgb[1015] = 24'b111011100100010000000000;
rgb[1016] = 24'b111111100101010100010001;
rgb[1017] = 24'b111111110110110100110010;
rgb[1018] = 24'b111111101000010101010101;
rgb[1019] = 24'b111111111001110101110110;
rgb[1020] = 24'b111111111011011010011001;
rgb[1021] = 24'b111111111100111010111011;
rgb[1022] = 24'b111111111110011011011101;
rgb[1023] = 24'b111111111111111111111111;
rgb[1024] = 24'b000000000000000000000000;
rgb[1025] = 24'b000100010001000100010001;
rgb[1026] = 24'b001000100010001000100010;
rgb[1027] = 24'b001100110011001100110011;
rgb[1028] = 24'b010001000100010001000100;
rgb[1029] = 24'b010101010101010101010101;
rgb[1030] = 24'b011001100110011001100110;
rgb[1031] = 24'b011101110111011101110111;
rgb[1032] = 24'b100010001000100010001000;
rgb[1033] = 24'b100110011001100110011001;
rgb[1034] = 24'b101010101010101010101010;
rgb[1035] = 24'b101110111011101110111011;
rgb[1036] = 24'b110011001100110011001100;
rgb[1037] = 24'b110111011101110111011101;
rgb[1038] = 24'b111011101110111011101110;
rgb[1039] = 24'b111111111111111111111111;
rgb[1040] = 24'b000000000000000000000000;
rgb[1041] = 24'b000100100001000000001111;
rgb[1042] = 24'b001001000010000100011111;
rgb[1043] = 24'b001101100011001000101111;
rgb[1044] = 24'b010010000100001000111111;
rgb[1045] = 24'b010110100101001101001111;
rgb[1046] = 24'b011011000110010001011111;
rgb[1047] = 24'b011111100111010101101111;
rgb[1048] = 24'b100011111000011010000000;
rgb[1049] = 24'b100111111001011110010010;
rgb[1050] = 24'b101011111010100010100100;
rgb[1051] = 24'b101111111011100110110110;
rgb[1052] = 24'b110011111100101111001000;
rgb[1053] = 24'b110111111101110011011010;
rgb[1054] = 24'b111011111110110111101100;
rgb[1055] = 24'b111111111111111111111111;
rgb[1056] = 24'b000000000000000000000000;
rgb[1057] = 24'b000100110001000000001110;
rgb[1058] = 24'b001001100010000000011101;
rgb[1059] = 24'b001110010011000100101100;
rgb[1060] = 24'b010011010100000100111010;
rgb[1061] = 24'b011000000101001001001001;
rgb[1062] = 24'b011100110110001001011000;
rgb[1063] = 24'b100001100111001101100111;
rgb[1064] = 24'b100101111000010001111000;
rgb[1065] = 24'b101001101001010110001011;
rgb[1066] = 24'b101101011010011110011110;
rgb[1067] = 24'b110001001011100010110001;
rgb[1068] = 24'b110100101100101011000101;
rgb[1069] = 24'b111000011101101111011000;
rgb[1070] = 24'b111100001110110111101011;
rgb[1071] = 24'b111111111111111111111111;
rgb[1072] = 24'b000000000000000000000000;
rgb[1073] = 24'b000101000001000000001101;
rgb[1074] = 24'b001010000010000000011011;
rgb[1075] = 24'b001111010011000000101000;
rgb[1076] = 24'b010100010100000000110110;
rgb[1077] = 24'b011001010101000001000100;
rgb[1078] = 24'b011110100110000101010001;
rgb[1079] = 24'b100011100111000101011111;
rgb[1080] = 24'b100111111000001001110000;
rgb[1081] = 24'b101011011001010010000100;
rgb[1082] = 24'b101110111010010110011000;
rgb[1083] = 24'b110010001011011110101101;
rgb[1084] = 24'b110101101100100111000001;
rgb[1085] = 24'b111000111101101111010110;
rgb[1086] = 24'b111100011110110111101010;
rgb[1087] = 24'b111111111111111111111111;
rgb[1088] = 24'b000000000000000000000000;
rgb[1089] = 24'b000101010000111100001100;
rgb[1090] = 24'b001010110001111100011000;
rgb[1091] = 24'b010000000010111100100101;
rgb[1092] = 24'b010101100011111100110001;
rgb[1093] = 24'b011010110100111100111110;
rgb[1094] = 24'b100000010101111101001010;
rgb[1095] = 24'b100101100110111101010111;
rgb[1096] = 24'b101001111000000001101000;
rgb[1097] = 24'b101101001001001001111101;
rgb[1098] = 24'b110000001010010010010011;
rgb[1099] = 24'b110011011011011010101000;
rgb[1100] = 24'b110110011100100010111110;
rgb[1101] = 24'b111001101101101011010011;
rgb[1102] = 24'b111100101110110011101001;
rgb[1103] = 24'b111111111111111111111111;
rgb[1104] = 24'b000000000000000000000000;
rgb[1105] = 24'b000101100000111100001011;
rgb[1106] = 24'b001011010001111100010110;
rgb[1107] = 24'b010001000010111000100010;
rgb[1108] = 24'b010110100011111000101101;
rgb[1109] = 24'b011100010100111000111000;
rgb[1110] = 24'b100010000101110101000100;
rgb[1111] = 24'b100111100110110101001111;
rgb[1112] = 24'b101011110111111001100000;
rgb[1113] = 24'b101110111001000001110110;
rgb[1114] = 24'b110001101010001110001101;
rgb[1115] = 24'b110100011011010110100100;
rgb[1116] = 24'b110111011100011110111011;
rgb[1117] = 24'b111010001101101011010001;
rgb[1118] = 24'b111100111110110011101000;
rgb[1119] = 24'b111111111111111111111111;
rgb[1120] = 24'b000000000000000000000000;
rgb[1121] = 24'b000101110000111100001010;
rgb[1122] = 24'b001011110001111000010100;
rgb[1123] = 24'b010001110010111000011110;
rgb[1124] = 24'b010111110011110100101000;
rgb[1125] = 24'b011101100100110000110011;
rgb[1126] = 24'b100011100101110000111101;
rgb[1127] = 24'b101001100110101101000111;
rgb[1128] = 24'b101101110111110001011000;
rgb[1129] = 24'b110000011000111101110000;
rgb[1130] = 24'b110011001010000110000111;
rgb[1131] = 24'b110101101011010010011111;
rgb[1132] = 24'b111000001100011110110111;
rgb[1133] = 24'b111010101101100111001111;
rgb[1134] = 24'b111101001110110011100111;
rgb[1135] = 24'b111111101111111111111111;
rgb[1136] = 24'b000000000000000000000000;
rgb[1137] = 24'b000110000000111100001001;
rgb[1138] = 24'b001100010001111000010010;
rgb[1139] = 24'b010010100010110100011011;
rgb[1140] = 24'b011000110011110000100100;
rgb[1141] = 24'b011111000100101100101101;
rgb[1142] = 24'b100101010101101000110110;
rgb[1143] = 24'b101011100110100100111111;
rgb[1144] = 24'b101111110111101001010000;
rgb[1145] = 24'b110010001000110101101001;
rgb[1146] = 24'b110100011010000010000010;
rgb[1147] = 24'b110110101011001110011011;
rgb[1148] = 24'b111000111100011010110100;
rgb[1149] = 24'b111011001101100111001101;
rgb[1150] = 24'b111101011110110011100110;
rgb[1151] = 24'b111111111111111111111111;
rgb[1152] = 24'b000000000000000000000000;
rgb[1153] = 24'b000110100000111000000111;
rgb[1154] = 24'b001101000001110100001111;
rgb[1155] = 24'b010011100010110000010111;
rgb[1156] = 24'b011010000011101100011111;
rgb[1157] = 24'b100000100100101000100111;
rgb[1158] = 24'b100111000101100100101111;
rgb[1159] = 24'b101101100110011100110111;
rgb[1160] = 24'b110001110111100001001000;
rgb[1161] = 24'b110011111000110001100010;
rgb[1162] = 24'b110101111001111101111100;
rgb[1163] = 24'b110111111011001010010110;
rgb[1164] = 24'b111001111100010110110000;
rgb[1165] = 24'b111011111101100011001010;
rgb[1166] = 24'b111101111110101111100100;
rgb[1167] = 24'b111111101111111111111111;
rgb[1168] = 24'b000000000000000000000000;
rgb[1169] = 24'b000110110000111000000110;
rgb[1170] = 24'b001101100001110100001101;
rgb[1171] = 24'b010100010010101100010100;
rgb[1172] = 24'b011011000011101000011011;
rgb[1173] = 24'b100010000100100000100001;
rgb[1174] = 24'b101000110101011100101000;
rgb[1175] = 24'b101111100110010100101111;
rgb[1176] = 24'b110011110111011101000000;
rgb[1177] = 24'b110101101000101001011011;
rgb[1178] = 24'b110111011001110101110110;
rgb[1179] = 24'b111000111011000110010010;
rgb[1180] = 24'b111010101100010010101101;
rgb[1181] = 24'b111100011101100011001000;
rgb[1182] = 24'b111110001110101111100011;
rgb[1183] = 24'b111111111111111111111111;
rgb[1184] = 24'b000000000000000000000000;
rgb[1185] = 24'b000111000000111000000101;
rgb[1186] = 24'b001110000001110000001011;
rgb[1187] = 24'b010101010010101000010001;
rgb[1188] = 24'b011100010011100100010110;
rgb[1189] = 24'b100011010100011100011100;
rgb[1190] = 24'b101010100101010100100010;
rgb[1191] = 24'b110001100110010000100111;
rgb[1192] = 24'b110101110111010100111000;
rgb[1193] = 24'b110111011000100001010100;
rgb[1194] = 24'b111000101001110001110001;
rgb[1195] = 24'b111010001011000010001101;
rgb[1196] = 24'b111011101100001110101010;
rgb[1197] = 24'b111100111101011111000110;
rgb[1198] = 24'b111110011110101111100010;
rgb[1199] = 24'b111111101111111111111111;
rgb[1200] = 24'b000000000000000000000000;
rgb[1201] = 24'b000111010000111000000100;
rgb[1202] = 24'b001110100001110000001001;
rgb[1203] = 24'b010110000010101000001101;
rgb[1204] = 24'b011101010011100000010010;
rgb[1205] = 24'b100100110100011000010110;
rgb[1206] = 24'b101100000101010000011011;
rgb[1207] = 24'b110011100110001000011111;
rgb[1208] = 24'b110111110111001100110000;
rgb[1209] = 24'b111000111000011101001110;
rgb[1210] = 24'b111010001001101101101011;
rgb[1211] = 24'b111011001010111110001001;
rgb[1212] = 24'b111100011100001110100110;
rgb[1213] = 24'b111101011101011111000100;
rgb[1214] = 24'b111110101110101111100001;
rgb[1215] = 24'b111111111111111111111111;
rgb[1216] = 24'b000000000000000000000000;
rgb[1217] = 24'b000111100000110100000011;
rgb[1218] = 24'b001111010001101100000110;
rgb[1219] = 24'b010110110010100100001010;
rgb[1220] = 24'b011110100011011100001101;
rgb[1221] = 24'b100110010100010000010000;
rgb[1222] = 24'b101101110101001000010100;
rgb[1223] = 24'b110101100110000000010111;
rgb[1224] = 24'b111001110111000100101000;
rgb[1225] = 24'b111010101000010101000111;
rgb[1226] = 24'b111011101001100101100101;
rgb[1227] = 24'b111100011010111010000100;
rgb[1228] = 24'b111101001100001010100011;
rgb[1229] = 24'b111110001101011011000001;
rgb[1230] = 24'b111110111110101011100000;
rgb[1231] = 24'b111111111111111111111111;
rgb[1232] = 24'b000000000000000000000000;
rgb[1233] = 24'b000111110000110100000010;
rgb[1234] = 24'b001111110001101000000100;
rgb[1235] = 24'b010111110010100000000110;
rgb[1236] = 24'b011111100011010100001001;
rgb[1237] = 24'b100111100100001100001011;
rgb[1238] = 24'b101111100101000000001101;
rgb[1239] = 24'b110111100101111000001111;
rgb[1240] = 24'b111011110110111100100000;
rgb[1241] = 24'b111100011000001101000000;
rgb[1242] = 24'b111100111001100001100000;
rgb[1243] = 24'b111101011010110010000000;
rgb[1244] = 24'b111110001100000110011111;
rgb[1245] = 24'b111110101101010110111111;
rgb[1246] = 24'b111111001110101011011111;
rgb[1247] = 24'b111111111111111111111111;
rgb[1248] = 24'b000000000000000000000000;
rgb[1249] = 24'b001000000000110100000001;
rgb[1250] = 24'b010000010001101000000010;
rgb[1251] = 24'b011000100010011100000011;
rgb[1252] = 24'b100000110011010000000100;
rgb[1253] = 24'b101001000100001000000101;
rgb[1254] = 24'b110001010100111100000110;
rgb[1255] = 24'b111001100101110000000111;
rgb[1256] = 24'b111101110110110100011000;
rgb[1257] = 24'b111110001000001000111001;
rgb[1258] = 24'b111110011001011101011010;
rgb[1259] = 24'b111110101010101101111011;
rgb[1260] = 24'b111110111100000010011100;
rgb[1261] = 24'b111111001101010110111101;
rgb[1262] = 24'b111111011110101011011110;
rgb[1263] = 24'b111111111111111111111111;
rgb[1264] = 24'b000000000000000000000000;
rgb[1265] = 24'b001000100000110000000000;
rgb[1266] = 24'b010001000001100100000000;
rgb[1267] = 24'b011001100010011000000000;
rgb[1268] = 24'b100010000011001100000000;
rgb[1269] = 24'b101010100100000000000000;
rgb[1270] = 24'b110011000100110100000000;
rgb[1271] = 24'b111011100101101000000000;
rgb[1272] = 24'b111111100110101100010001;
rgb[1273] = 24'b111111111000000000110010;
rgb[1274] = 24'b111111101001010101010101;
rgb[1275] = 24'b111111111010101001110110;
rgb[1276] = 24'b111111111011111110011001;
rgb[1277] = 24'b111111111101010010111011;
rgb[1278] = 24'b111111111110100111011101;
rgb[1279] = 24'b111111111111111111111111;
rgb[1280] = 24'b000000000000000000000000;
rgb[1281] = 24'b000100010001000100010001;
rgb[1282] = 24'b001000100010001000100010;
rgb[1283] = 24'b001100110011001100110011;
rgb[1284] = 24'b010001000100010001000100;
rgb[1285] = 24'b010101010101010101010101;
rgb[1286] = 24'b011001100110011001100110;
rgb[1287] = 24'b011101110111011101110111;
rgb[1288] = 24'b100010001000100010001000;
rgb[1289] = 24'b100110011001100110011001;
rgb[1290] = 24'b101010101010101010101010;
rgb[1291] = 24'b101110111011101110111011;
rgb[1292] = 24'b110011001100110011001100;
rgb[1293] = 24'b110111011101110111011101;
rgb[1294] = 24'b111011101110111011101110;
rgb[1295] = 24'b111111111111111111111111;
rgb[1296] = 24'b000000000000000000000000;
rgb[1297] = 24'b000100100001000000001111;
rgb[1298] = 24'b001001000010000100011111;
rgb[1299] = 24'b001101100011001000101111;
rgb[1300] = 24'b010010000100001100111111;
rgb[1301] = 24'b010110100101010001001111;
rgb[1302] = 24'b011011000110010101011111;
rgb[1303] = 24'b011111100111011001101111;
rgb[1304] = 24'b100011111000011110000000;
rgb[1305] = 24'b100111111001100010010010;
rgb[1306] = 24'b101011111010100110100100;
rgb[1307] = 24'b101111111011101010110110;
rgb[1308] = 24'b110011111100101111001000;
rgb[1309] = 24'b110111111101110011011010;
rgb[1310] = 24'b111011111110110111101100;
rgb[1311] = 24'b111111111111111111111111;
rgb[1312] = 24'b000000000000000000000000;
rgb[1313] = 24'b000100110001000000001110;
rgb[1314] = 24'b001001100010000100011101;
rgb[1315] = 24'b001110010011001000101100;
rgb[1316] = 24'b010011010100001100111010;
rgb[1317] = 24'b011000000101010001001001;
rgb[1318] = 24'b011100110110010101011000;
rgb[1319] = 24'b100001100111011001100111;
rgb[1320] = 24'b100101111000011101111000;
rgb[1321] = 24'b101001101001100010001011;
rgb[1322] = 24'b101101011010100110011110;
rgb[1323] = 24'b110001001011101010110001;
rgb[1324] = 24'b110100101100101111000101;
rgb[1325] = 24'b111000011101110011011000;
rgb[1326] = 24'b111100001110110111101011;
rgb[1327] = 24'b111111111111111111111111;
rgb[1328] = 24'b000000000000000000000000;
rgb[1329] = 24'b000101000001000000001101;
rgb[1330] = 24'b001010000010000100011011;
rgb[1331] = 24'b001111010011001000101000;
rgb[1332] = 24'b010100010100001100110110;
rgb[1333] = 24'b011001010101010001000100;
rgb[1334] = 24'b011110100110010101010001;
rgb[1335] = 24'b100011100111010101011111;
rgb[1336] = 24'b100111111000011001110000;
rgb[1337] = 24'b101011011001100010000100;
rgb[1338] = 24'b101110111010100110011000;
rgb[1339] = 24'b110010001011101010101101;
rgb[1340] = 24'b110101101100101111000001;
rgb[1341] = 24'b111000111101110011010110;
rgb[1342] = 24'b111100011110110111101010;
rgb[1343] = 24'b111111111111111111111111;
rgb[1344] = 24'b000000000000000000000000;
rgb[1345] = 24'b000101010001000000001100;
rgb[1346] = 24'b001010110010000100011000;
rgb[1347] = 24'b010000000011001000100101;
rgb[1348] = 24'b010101100100001100110001;
rgb[1349] = 24'b011010110101001100111110;
rgb[1350] = 24'b100000010110010001001010;
rgb[1351] = 24'b100101100111010101010111;
rgb[1352] = 24'b101001111000011001101000;
rgb[1353] = 24'b101101001001011101111101;
rgb[1354] = 24'b110000001010100010010011;
rgb[1355] = 24'b110011011011101010101000;
rgb[1356] = 24'b110110011100101110111110;
rgb[1357] = 24'b111001101101110011010011;
rgb[1358] = 24'b111100101110110111101001;
rgb[1359] = 24'b111111111111111111111111;
rgb[1360] = 24'b000000000000000000000000;
rgb[1361] = 24'b000101100001000000001011;
rgb[1362] = 24'b001011010010000100010110;
rgb[1363] = 24'b010001000011001000100010;
rgb[1364] = 24'b010110100100001000101101;
rgb[1365] = 24'b011100010101001100111000;
rgb[1366] = 24'b100010000110010001000100;
rgb[1367] = 24'b100111100111010101001111;
rgb[1368] = 24'b101011111000011001100000;
rgb[1369] = 24'b101110111001011101110110;
rgb[1370] = 24'b110001101010100010001101;
rgb[1371] = 24'b110100011011100110100100;
rgb[1372] = 24'b110111011100101110111011;
rgb[1373] = 24'b111010001101110011010001;
rgb[1374] = 24'b111100111110110111101000;
rgb[1375] = 24'b111111111111111111111111;
rgb[1376] = 24'b000000000000000000000000;
rgb[1377] = 24'b000101110001000000001010;
rgb[1378] = 24'b001011110010000100010100;
rgb[1379] = 24'b010001110011001000011110;
rgb[1380] = 24'b010111110100001000101000;
rgb[1381] = 24'b011101100101001100110011;
rgb[1382] = 24'b100011100110010000111101;
rgb[1383] = 24'b101001100111010001000111;
rgb[1384] = 24'b101101111000010101011000;
rgb[1385] = 24'b110000011001011101110000;
rgb[1386] = 24'b110011001010100010000111;
rgb[1387] = 24'b110101101011100110011111;
rgb[1388] = 24'b111000001100101110110111;
rgb[1389] = 24'b111010101101110011001111;
rgb[1390] = 24'b111101001110110111100111;
rgb[1391] = 24'b111111101111111111111111;
rgb[1392] = 24'b000000000000000000000000;
rgb[1393] = 24'b000110000001000000001001;
rgb[1394] = 24'b001100010010000100010010;
rgb[1395] = 24'b010010100011000100011011;
rgb[1396] = 24'b011000110100001000100100;
rgb[1397] = 24'b011111000101001100101101;
rgb[1398] = 24'b100101010110001100110110;
rgb[1399] = 24'b101011100111010000111111;
rgb[1400] = 24'b101111111000010101010000;
rgb[1401] = 24'b110010001001011001101001;
rgb[1402] = 24'b110100011010100010000010;
rgb[1403] = 24'b110110101011100110011011;
rgb[1404] = 24'b111000111100101010110100;
rgb[1405] = 24'b111011001101110011001101;
rgb[1406] = 24'b111101011110110111100110;
rgb[1407] = 24'b111111111111111111111111;
rgb[1408] = 24'b000000000000000000000000;
rgb[1409] = 24'b000110100001000000000111;
rgb[1410] = 24'b001101000010000100001111;
rgb[1411] = 24'b010011100011000100010111;
rgb[1412] = 24'b011010000100001000011111;
rgb[1413] = 24'b100000100101001000100111;
rgb[1414] = 24'b100111000110001100101111;
rgb[1415] = 24'b101101100111001100110111;
rgb[1416] = 24'b110001111000010001001000;
rgb[1417] = 24'b110011111001011001100010;
rgb[1418] = 24'b110101111010011101111100;
rgb[1419] = 24'b110111111011100110010110;
rgb[1420] = 24'b111001111100101010110000;
rgb[1421] = 24'b111011111101110011001010;
rgb[1422] = 24'b111101111110110111100100;
rgb[1423] = 24'b111111101111111111111111;
rgb[1424] = 24'b000000000000000000000000;
rgb[1425] = 24'b000110110001000000000110;
rgb[1426] = 24'b001101100010000100001101;
rgb[1427] = 24'b010100010011000100010100;
rgb[1428] = 24'b011011000100001000011011;
rgb[1429] = 24'b100010000101001000100001;
rgb[1430] = 24'b101000110110001100101000;
rgb[1431] = 24'b101111100111001100101111;
rgb[1432] = 24'b110011111000010001000000;
rgb[1433] = 24'b110101101001011001011011;
rgb[1434] = 24'b110111011010011101110110;
rgb[1435] = 24'b111000111011100110010010;
rgb[1436] = 24'b111010101100101010101101;
rgb[1437] = 24'b111100011101110011001000;
rgb[1438] = 24'b111110001110110111100011;
rgb[1439] = 24'b111111111111111111111111;
rgb[1440] = 24'b000000000000000000000000;
rgb[1441] = 24'b000111000001000000000101;
rgb[1442] = 24'b001110000010000000001011;
rgb[1443] = 24'b010101010011000100010001;
rgb[1444] = 24'b011100010100000100010110;
rgb[1445] = 24'b100011010101001000011100;
rgb[1446] = 24'b101010100110001000100010;
rgb[1447] = 24'b110001100111001100100111;
rgb[1448] = 24'b110101111000010000111000;
rgb[1449] = 24'b110111011001010101010100;
rgb[1450] = 24'b111000101010011101110001;
rgb[1451] = 24'b111010001011100010001101;
rgb[1452] = 24'b111011101100101010101010;
rgb[1453] = 24'b111100111101101111000110;
rgb[1454] = 24'b111110011110110111100010;
rgb[1455] = 24'b111111101111111111111111;
rgb[1456] = 24'b000000000000000000000000;
rgb[1457] = 24'b000111010001000000000100;
rgb[1458] = 24'b001110100010000000001001;
rgb[1459] = 24'b010110000011000100001101;
rgb[1460] = 24'b011101010100000100010010;
rgb[1461] = 24'b100100110101001000010110;
rgb[1462] = 24'b101100000110001000011011;
rgb[1463] = 24'b110011100111001000011111;
rgb[1464] = 24'b110111111000001100110000;
rgb[1465] = 24'b111000111001010101001110;
rgb[1466] = 24'b111010001010011101101011;
rgb[1467] = 24'b111011001011100010001001;
rgb[1468] = 24'b111100011100101010100110;
rgb[1469] = 24'b111101011101101111000100;
rgb[1470] = 24'b111110101110110111100001;
rgb[1471] = 24'b111111111111111111111111;
rgb[1472] = 24'b000000000000000000000000;
rgb[1473] = 24'b000111100001000000000011;
rgb[1474] = 24'b001111010010000000000110;
rgb[1475] = 24'b010110110011000100001010;
rgb[1476] = 24'b011110100100000100001101;
rgb[1477] = 24'b100110010101000100010000;
rgb[1478] = 24'b101101110110001000010100;
rgb[1479] = 24'b110101100111001000010111;
rgb[1480] = 24'b111001111000001100101000;
rgb[1481] = 24'b111010101001010101000111;
rgb[1482] = 24'b111011101010011001100101;
rgb[1483] = 24'b111100011011100010000100;
rgb[1484] = 24'b111101001100101010100011;
rgb[1485] = 24'b111110001101101111000001;
rgb[1486] = 24'b111110111110110111100000;
rgb[1487] = 24'b111111111111111111111111;
rgb[1488] = 24'b000000000000000000000000;
rgb[1489] = 24'b000111110001000000000010;
rgb[1490] = 24'b001111110010000000000100;
rgb[1491] = 24'b010111110011000000000110;
rgb[1492] = 24'b011111100100000100001001;
rgb[1493] = 24'b100111100101000100001011;
rgb[1494] = 24'b101111100110000100001101;
rgb[1495] = 24'b110111100111001000001111;
rgb[1496] = 24'b111011111000001100100000;
rgb[1497] = 24'b111100011001010001000000;
rgb[1498] = 24'b111100111010011001100000;
rgb[1499] = 24'b111101011011100010000000;
rgb[1500] = 24'b111110001100100110011111;
rgb[1501] = 24'b111110101101101110111111;
rgb[1502] = 24'b111111001110110111011111;
rgb[1503] = 24'b111111111111111111111111;
rgb[1504] = 24'b000000000000000000000000;
rgb[1505] = 24'b001000000001000000000001;
rgb[1506] = 24'b010000010010000000000010;
rgb[1507] = 24'b011000100011000000000011;
rgb[1508] = 24'b100000110100000000000100;
rgb[1509] = 24'b101001000101000100000101;
rgb[1510] = 24'b110001010110000100000110;
rgb[1511] = 24'b111001100111000100000111;
rgb[1512] = 24'b111101111000001000011000;
rgb[1513] = 24'b111110001001010000111001;
rgb[1514] = 24'b111110011010011001011010;
rgb[1515] = 24'b111110101011011101111011;
rgb[1516] = 24'b111110111100100110011100;
rgb[1517] = 24'b111111001101101110111101;
rgb[1518] = 24'b111111011110110111011110;
rgb[1519] = 24'b111111111111111111111111;
rgb[1520] = 24'b000000000000000000000000;
rgb[1521] = 24'b001000100001000000000000;
rgb[1522] = 24'b010001000010000000000000;
rgb[1523] = 24'b011001100011000000000000;
rgb[1524] = 24'b100010000100000000000000;
rgb[1525] = 24'b101010100101000000000000;
rgb[1526] = 24'b110011000110000100000000;
rgb[1527] = 24'b111011100111000100000000;
rgb[1528] = 24'b111111101000001000010001;
rgb[1529] = 24'b111111111001010000110010;
rgb[1530] = 24'b111111101010010101010101;
rgb[1531] = 24'b111111111011011101110110;
rgb[1532] = 24'b111111111100100110011001;
rgb[1533] = 24'b111111111101101110111011;
rgb[1534] = 24'b111111111110110111011101;
rgb[1535] = 24'b111111111111111111111111;
rgb[1536] = 24'b000000000000000000000000;
rgb[1537] = 24'b000100010001000100010001;
rgb[1538] = 24'b001000100010001000100010;
rgb[1539] = 24'b001100110011001100110011;
rgb[1540] = 24'b010001000100010001000100;
rgb[1541] = 24'b010101010101010101010101;
rgb[1542] = 24'b011001100110011001100110;
rgb[1543] = 24'b011101110111011101110111;
rgb[1544] = 24'b100010001000100010001000;
rgb[1545] = 24'b100110011001100110011001;
rgb[1546] = 24'b101010101010101010101010;
rgb[1547] = 24'b101110111011101110111011;
rgb[1548] = 24'b110011001100110011001100;
rgb[1549] = 24'b110111011101110111011101;
rgb[1550] = 24'b111011101110111011101110;
rgb[1551] = 24'b111111111111111111111111;
rgb[1552] = 24'b000000000000000000000000;
rgb[1553] = 24'b000100100001000100001111;
rgb[1554] = 24'b001001000010001000011111;
rgb[1555] = 24'b001101100011001100101111;
rgb[1556] = 24'b010010000100010000111111;
rgb[1557] = 24'b010110100101010101001111;
rgb[1558] = 24'b011011000110011001011111;
rgb[1559] = 24'b011111100111100001101111;
rgb[1560] = 24'b100011111000100110000000;
rgb[1561] = 24'b100111111001100110010010;
rgb[1562] = 24'b101011111010101010100100;
rgb[1563] = 24'b101111111011101110110110;
rgb[1564] = 24'b110011111100110011001000;
rgb[1565] = 24'b110111111101110111011010;
rgb[1566] = 24'b111011111110111011101100;
rgb[1567] = 24'b111111111111111111111111;
rgb[1568] = 24'b000000000000000000000000;
rgb[1569] = 24'b000100110001000100001110;
rgb[1570] = 24'b001001100010001000011101;
rgb[1571] = 24'b001110010011001100101100;
rgb[1572] = 24'b010011010100010100111010;
rgb[1573] = 24'b011000000101011001001001;
rgb[1574] = 24'b011100110110011101011000;
rgb[1575] = 24'b100001100111100101100111;
rgb[1576] = 24'b100101111000101001111000;
rgb[1577] = 24'b101001101001101010001011;
rgb[1578] = 24'b101101011010101110011110;
rgb[1579] = 24'b110001001011110010110001;
rgb[1580] = 24'b110100101100110011000101;
rgb[1581] = 24'b111000011101110111011000;
rgb[1582] = 24'b111100001110111011101011;
rgb[1583] = 24'b111111111111111111111111;
rgb[1584] = 24'b000000000000000000000000;
rgb[1585] = 24'b000101000001000100001101;
rgb[1586] = 24'b001010000010001000011011;
rgb[1587] = 24'b001111010011010000101000;
rgb[1588] = 24'b010100010100010100110110;
rgb[1589] = 24'b011001010101011101000100;
rgb[1590] = 24'b011110100110100001010001;
rgb[1591] = 24'b100011100111101001011111;
rgb[1592] = 24'b100111111000101101110000;
rgb[1593] = 24'b101011011001101110000100;
rgb[1594] = 24'b101110111010110010011000;
rgb[1595] = 24'b110010001011110010101101;
rgb[1596] = 24'b110101101100110111000001;
rgb[1597] = 24'b111000111101110111010110;
rgb[1598] = 24'b111100011110111011101010;
rgb[1599] = 24'b111111111111111111111111;
rgb[1600] = 24'b000000000000000000000000;
rgb[1601] = 24'b000101010001000100001100;
rgb[1602] = 24'b001010110010001100011000;
rgb[1603] = 24'b010000000011010000100101;
rgb[1604] = 24'b010101100100011000110001;
rgb[1605] = 24'b011010110101100000111110;
rgb[1606] = 24'b100000010110100101001010;
rgb[1607] = 24'b100101100111101101010111;
rgb[1608] = 24'b101001111000110001101000;
rgb[1609] = 24'b101101001001110001111101;
rgb[1610] = 24'b110000001010110110010011;
rgb[1611] = 24'b110011011011110110101000;
rgb[1612] = 24'b110110011100110110111110;
rgb[1613] = 24'b111001101101111011010011;
rgb[1614] = 24'b111100101110111011101001;
rgb[1615] = 24'b111111111111111111111111;
rgb[1616] = 24'b000000000000000000000000;
rgb[1617] = 24'b000101100001000100001011;
rgb[1618] = 24'b001011010010001100010110;
rgb[1619] = 24'b010001000011010100100010;
rgb[1620] = 24'b010110100100011100101101;
rgb[1621] = 24'b011100010101100100111000;
rgb[1622] = 24'b100010000110101001000100;
rgb[1623] = 24'b100111100111110001001111;
rgb[1624] = 24'b101011111000110101100000;
rgb[1625] = 24'b101110111001110101110110;
rgb[1626] = 24'b110001101010111010001101;
rgb[1627] = 24'b110100011011111010100100;
rgb[1628] = 24'b110111011100111010111011;
rgb[1629] = 24'b111010001101111011010001;
rgb[1630] = 24'b111100111110111011101000;
rgb[1631] = 24'b111111111111111111111111;
rgb[1632] = 24'b000000000000000000000000;
rgb[1633] = 24'b000101110001000100001010;
rgb[1634] = 24'b001011110010001100010100;
rgb[1635] = 24'b010001110011010100011110;
rgb[1636] = 24'b010111110100011100101000;
rgb[1637] = 24'b011101100101100100110011;
rgb[1638] = 24'b100011100110101100111101;
rgb[1639] = 24'b101001100111110101000111;
rgb[1640] = 24'b101101111000111001011000;
rgb[1641] = 24'b110000011001111001110000;
rgb[1642] = 24'b110011001010111010000111;
rgb[1643] = 24'b110101101011111010011111;
rgb[1644] = 24'b111000001100111010110111;
rgb[1645] = 24'b111010101101111011001111;
rgb[1646] = 24'b111101001110111011100111;
rgb[1647] = 24'b111111101111111011111111;
rgb[1648] = 24'b000000000000000000000000;
rgb[1649] = 24'b000110000001001000001001;
rgb[1650] = 24'b001100010010010000010010;
rgb[1651] = 24'b010010100011011000011011;
rgb[1652] = 24'b011000110100100000100100;
rgb[1653] = 24'b011111000101101000101101;
rgb[1654] = 24'b100101010110110000110110;
rgb[1655] = 24'b101011100111111000111111;
rgb[1656] = 24'b101111111000111101010000;
rgb[1657] = 24'b110010001001111101101001;
rgb[1658] = 24'b110100011010111110000010;
rgb[1659] = 24'b110110101011111110011011;
rgb[1660] = 24'b111000111100111110110100;
rgb[1661] = 24'b111011001101111111001101;
rgb[1662] = 24'b111101011110111111100110;
rgb[1663] = 24'b111111111111111111111111;
rgb[1664] = 24'b000000000000000000000000;
rgb[1665] = 24'b000110100001001000000111;
rgb[1666] = 24'b001101000010010000001111;
rgb[1667] = 24'b010011100011011000010111;
rgb[1668] = 24'b011010000100100100011111;
rgb[1669] = 24'b100000100101101100100111;
rgb[1670] = 24'b100111000110110100101111;
rgb[1671] = 24'b101101101000000000110111;
rgb[1672] = 24'b110001111001000101001000;
rgb[1673] = 24'b110011111010000001100010;
rgb[1674] = 24'b110101111011000001111100;
rgb[1675] = 24'b110111111100000010010110;
rgb[1676] = 24'b111001111100111110110000;
rgb[1677] = 24'b111011111101111111001010;
rgb[1678] = 24'b111101111110111111100100;
rgb[1679] = 24'b111111101111111011111111;
rgb[1680] = 24'b000000000000000000000000;
rgb[1681] = 24'b000110110001001000000110;
rgb[1682] = 24'b001101100010010000001101;
rgb[1683] = 24'b010100010011011100010100;
rgb[1684] = 24'b011011000100100100011011;
rgb[1685] = 24'b100010000101110000100001;
rgb[1686] = 24'b101000110110111000101000;
rgb[1687] = 24'b101111101000000100101111;
rgb[1688] = 24'b110011111001001001000000;
rgb[1689] = 24'b110101101010000101011011;
rgb[1690] = 24'b110111011011000101110110;
rgb[1691] = 24'b111000111100000010010010;
rgb[1692] = 24'b111010101101000010101101;
rgb[1693] = 24'b111100011101111111001000;
rgb[1694] = 24'b111110001110111111100011;
rgb[1695] = 24'b111111111111111111111111;
rgb[1696] = 24'b000000000000000000000000;
rgb[1697] = 24'b000111000001001000000101;
rgb[1698] = 24'b001110000010010100001011;
rgb[1699] = 24'b010101010011011100010001;
rgb[1700] = 24'b011100010100101000010110;
rgb[1701] = 24'b100011010101110100011100;
rgb[1702] = 24'b101010100110111100100010;
rgb[1703] = 24'b110001101000001000100111;
rgb[1704] = 24'b110101111001001100111000;
rgb[1705] = 24'b110111011010001001010100;
rgb[1706] = 24'b111000101011001001110001;
rgb[1707] = 24'b111010001100000110001101;
rgb[1708] = 24'b111011101101000010101010;
rgb[1709] = 24'b111100111110000011000110;
rgb[1710] = 24'b111110011110111111100010;
rgb[1711] = 24'b111111101111111011111111;
rgb[1712] = 24'b000000000000000000000000;
rgb[1713] = 24'b000111010001001000000100;
rgb[1714] = 24'b001110100010010100001001;
rgb[1715] = 24'b010110000011100000001101;
rgb[1716] = 24'b011101010100101100010010;
rgb[1717] = 24'b100100110101110100010110;
rgb[1718] = 24'b101100000111000000011011;
rgb[1719] = 24'b110011101000001100011111;
rgb[1720] = 24'b110111111001010000110000;
rgb[1721] = 24'b111000111010001101001110;
rgb[1722] = 24'b111010001011001001101011;
rgb[1723] = 24'b111011001100001010001001;
rgb[1724] = 24'b111100011101000110100110;
rgb[1725] = 24'b111101011110000011000100;
rgb[1726] = 24'b111110101110111111100001;
rgb[1727] = 24'b111111111111111111111111;
rgb[1728] = 24'b000000000000000000000000;
rgb[1729] = 24'b000111100001001000000011;
rgb[1730] = 24'b001111010010010100000110;
rgb[1731] = 24'b010110110011100000001010;
rgb[1732] = 24'b011110100100101100001101;
rgb[1733] = 24'b100110010101111000010000;
rgb[1734] = 24'b101101110111000100010100;
rgb[1735] = 24'b110101101000010000010111;
rgb[1736] = 24'b111001111001010100101000;
rgb[1737] = 24'b111010101010010001000111;
rgb[1738] = 24'b111011101011001101100101;
rgb[1739] = 24'b111100011100001010000100;
rgb[1740] = 24'b111101001101000110100011;
rgb[1741] = 24'b111110001110000011000001;
rgb[1742] = 24'b111110111110111111100000;
rgb[1743] = 24'b111111111111111111111111;
rgb[1744] = 24'b000000000000000000000000;
rgb[1745] = 24'b000111110001001100000010;
rgb[1746] = 24'b001111110010011000000100;
rgb[1747] = 24'b010111110011100100000110;
rgb[1748] = 24'b011111100100110000001001;
rgb[1749] = 24'b100111100101111100001011;
rgb[1750] = 24'b101111100111001000001101;
rgb[1751] = 24'b110111101000010100001111;
rgb[1752] = 24'b111011111001011000100000;
rgb[1753] = 24'b111100011010010101000000;
rgb[1754] = 24'b111100111011010001100000;
rgb[1755] = 24'b111101011100001110000000;
rgb[1756] = 24'b111110001101001010011111;
rgb[1757] = 24'b111110101110000110111111;
rgb[1758] = 24'b111111001111000011011111;
rgb[1759] = 24'b111111111111111111111111;
rgb[1760] = 24'b000000000000000000000000;
rgb[1761] = 24'b001000000001001100000001;
rgb[1762] = 24'b010000010010011000000010;
rgb[1763] = 24'b011000100011100100000011;
rgb[1764] = 24'b100000110100110100000100;
rgb[1765] = 24'b101001000110000000000101;
rgb[1766] = 24'b110001010111001100000110;
rgb[1767] = 24'b111001101000011000000111;
rgb[1768] = 24'b111101111001011100011000;
rgb[1769] = 24'b111110001010011000111001;
rgb[1770] = 24'b111110011011010101011010;
rgb[1771] = 24'b111110101100010001111011;
rgb[1772] = 24'b111110111101001010011100;
rgb[1773] = 24'b111111001110000110111101;
rgb[1774] = 24'b111111011111000011011110;
rgb[1775] = 24'b111111111111111111111111;
rgb[1776] = 24'b000000000000000000000000;
rgb[1777] = 24'b001000100001001100000000;
rgb[1778] = 24'b010001000010011000000000;
rgb[1779] = 24'b011001100011101000000000;
rgb[1780] = 24'b100010000100110100000000;
rgb[1781] = 24'b101010100110000100000000;
rgb[1782] = 24'b110011000111010000000000;
rgb[1783] = 24'b111011101000100000000000;
rgb[1784] = 24'b111111101001100100010001;
rgb[1785] = 24'b111111111010011100110010;
rgb[1786] = 24'b111111101011011001010101;
rgb[1787] = 24'b111111111100010001110110;
rgb[1788] = 24'b111111111101001110011001;
rgb[1789] = 24'b111111111110000110111011;
rgb[1790] = 24'b111111111111000011011101;
rgb[1791] = 24'b111111111111111111111111;
rgb[1792] = 24'b000000000000000000000000;
rgb[1793] = 24'b000100010001000100010001;
rgb[1794] = 24'b001000100010001000100010;
rgb[1795] = 24'b001100110011001100110011;
rgb[1796] = 24'b010001000100010001000100;
rgb[1797] = 24'b010101010101010101010101;
rgb[1798] = 24'b011001100110011001100110;
rgb[1799] = 24'b011101110111011101110111;
rgb[1800] = 24'b100010001000100010001000;
rgb[1801] = 24'b100110011001100110011001;
rgb[1802] = 24'b101010101010101010101010;
rgb[1803] = 24'b101110111011101110111011;
rgb[1804] = 24'b110011001100110011001100;
rgb[1805] = 24'b110111011101110111011101;
rgb[1806] = 24'b111011101110111011101110;
rgb[1807] = 24'b111111111111111111111111;
rgb[1808] = 24'b000000000000000000000000;
rgb[1809] = 24'b000100100001000100001111;
rgb[1810] = 24'b001001000010001000011111;
rgb[1811] = 24'b001101100011010000101111;
rgb[1812] = 24'b010010000100010100111111;
rgb[1813] = 24'b010110100101011001001111;
rgb[1814] = 24'b011011000110100001011111;
rgb[1815] = 24'b011111100111100101101111;
rgb[1816] = 24'b100011111000101010000000;
rgb[1817] = 24'b100111111001101110010010;
rgb[1818] = 24'b101011111010101110100100;
rgb[1819] = 24'b101111111011110010110110;
rgb[1820] = 24'b110011111100110111001000;
rgb[1821] = 24'b110111111101110111011010;
rgb[1822] = 24'b111011111110111011101100;
rgb[1823] = 24'b111111111111111111111111;
rgb[1824] = 24'b000000000000000000000000;
rgb[1825] = 24'b000100110001000100001110;
rgb[1826] = 24'b001001100010001100011101;
rgb[1827] = 24'b001110010011010100101100;
rgb[1828] = 24'b010011010100011100111010;
rgb[1829] = 24'b011000000101100001001001;
rgb[1830] = 24'b011100110110101001011000;
rgb[1831] = 24'b100001100111110001100111;
rgb[1832] = 24'b100101111000110101111000;
rgb[1833] = 24'b101001101001110110001011;
rgb[1834] = 24'b101101011010110110011110;
rgb[1835] = 24'b110001001011111010110001;
rgb[1836] = 24'b110100101100111011000101;
rgb[1837] = 24'b111000011101111011011000;
rgb[1838] = 24'b111100001110111011101011;
rgb[1839] = 24'b111111111111111111111111;
rgb[1840] = 24'b000000000000000000000000;
rgb[1841] = 24'b000101000001001000001101;
rgb[1842] = 24'b001010000010010000011011;
rgb[1843] = 24'b001111010011011000101000;
rgb[1844] = 24'b010100010100100000110110;
rgb[1845] = 24'b011001010101101001000100;
rgb[1846] = 24'b011110100110110001010001;
rgb[1847] = 24'b100011100111111001011111;
rgb[1848] = 24'b100111111000111101110000;
rgb[1849] = 24'b101011011001111110000100;
rgb[1850] = 24'b101110111010111110011000;
rgb[1851] = 24'b110010001011111110101101;
rgb[1852] = 24'b110101101100111111000001;
rgb[1853] = 24'b111000111101111111010110;
rgb[1854] = 24'b111100011110111111101010;
rgb[1855] = 24'b111111111111111111111111;
rgb[1856] = 24'b000000000000000000000000;
rgb[1857] = 24'b000101010001001000001100;
rgb[1858] = 24'b001010110010010100011000;
rgb[1859] = 24'b010000000011011100100101;
rgb[1860] = 24'b010101100100101000110001;
rgb[1861] = 24'b011010110101110000111110;
rgb[1862] = 24'b100000010110111101001010;
rgb[1863] = 24'b100101101000000101010111;
rgb[1864] = 24'b101001111001001001101000;
rgb[1865] = 24'b101101001010001001111101;
rgb[1866] = 24'b110000001011000110010011;
rgb[1867] = 24'b110011011100000110101000;
rgb[1868] = 24'b110110011101000010111110;
rgb[1869] = 24'b111001101110000011010011;
rgb[1870] = 24'b111100101110111111101001;
rgb[1871] = 24'b111111111111111111111111;
rgb[1872] = 24'b000000000000000000000000;
rgb[1873] = 24'b000101100001001000001011;
rgb[1874] = 24'b001011010010010100010110;
rgb[1875] = 24'b010001000011100000100010;
rgb[1876] = 24'b010110100100101100101101;
rgb[1877] = 24'b011100010101111000111000;
rgb[1878] = 24'b100010000111000101000100;
rgb[1879] = 24'b100111101000010001001111;
rgb[1880] = 24'b101011111001010101100000;
rgb[1881] = 24'b101110111010010001110110;
rgb[1882] = 24'b110001101011001110001101;
rgb[1883] = 24'b110100011100001010100100;
rgb[1884] = 24'b110111011101000110111011;
rgb[1885] = 24'b111010001110000011010001;
rgb[1886] = 24'b111100111110111111101000;
rgb[1887] = 24'b111111111111111111111111;
rgb[1888] = 24'b000000000000000000000000;
rgb[1889] = 24'b000101110001001100001010;
rgb[1890] = 24'b001011110010011000010100;
rgb[1891] = 24'b010001110011100100011110;
rgb[1892] = 24'b010111110100110100101000;
rgb[1893] = 24'b011101100110000000110011;
rgb[1894] = 24'b100011100111001100111101;
rgb[1895] = 24'b101001101000011001000111;
rgb[1896] = 24'b101101111001011101011000;
rgb[1897] = 24'b110000011010011001110000;
rgb[1898] = 24'b110011001011010110000111;
rgb[1899] = 24'b110101101100010010011111;
rgb[1900] = 24'b111000001101001010110111;
rgb[1901] = 24'b111010101110000111001111;
rgb[1902] = 24'b111101001111000011100111;
rgb[1903] = 24'b111111101111111011111111;
rgb[1904] = 24'b000000000000000000000000;
rgb[1905] = 24'b000110000001001100001001;
rgb[1906] = 24'b001100010010011100010010;
rgb[1907] = 24'b010010100011101000011011;
rgb[1908] = 24'b011000110100111000100100;
rgb[1909] = 24'b011111000110001000101101;
rgb[1910] = 24'b100101010111010100110110;
rgb[1911] = 24'b101011101000100100111111;
rgb[1912] = 24'b101111111001101001010000;
rgb[1913] = 24'b110010001010100001101001;
rgb[1914] = 24'b110100011011011110000010;
rgb[1915] = 24'b110110101100010110011011;
rgb[1916] = 24'b111000111101001110110100;
rgb[1917] = 24'b111011001110001011001101;
rgb[1918] = 24'b111101011111000011100110;
rgb[1919] = 24'b111111111111111111111111;
rgb[1920] = 24'b000000000000000000000000;
rgb[1921] = 24'b000110100001010000000111;
rgb[1922] = 24'b001101000010100000001111;
rgb[1923] = 24'b010011100011110000010111;
rgb[1924] = 24'b011010000101000000011111;
rgb[1925] = 24'b100000100110010000100111;
rgb[1926] = 24'b100111000111100000101111;
rgb[1927] = 24'b101101101000110000110111;
rgb[1928] = 24'b110001111001110101001000;
rgb[1929] = 24'b110011111010101101100010;
rgb[1930] = 24'b110101111011100101111100;
rgb[1931] = 24'b110111111100011110010110;
rgb[1932] = 24'b111001111101010110110000;
rgb[1933] = 24'b111011111110001111001010;
rgb[1934] = 24'b111101111111000111100100;
rgb[1935] = 24'b111111101111111011111111;
rgb[1936] = 24'b000000000000000000000000;
rgb[1937] = 24'b000110110001010000000110;
rgb[1938] = 24'b001101100010100000001101;
rgb[1939] = 24'b010100010011110100010100;
rgb[1940] = 24'b011011000101000100011011;
rgb[1941] = 24'b100010000110010100100001;
rgb[1942] = 24'b101000110111101000101000;
rgb[1943] = 24'b101111101000111000101111;
rgb[1944] = 24'b110011111001111101000000;
rgb[1945] = 24'b110101101010110101011011;
rgb[1946] = 24'b110111011011101101110110;
rgb[1947] = 24'b111000111100100010010010;
rgb[1948] = 24'b111010101101011010101101;
rgb[1949] = 24'b111100011110001111001000;
rgb[1950] = 24'b111110001111000111100011;
rgb[1951] = 24'b111111111111111111111111;
rgb[1952] = 24'b000000000000000000000000;
rgb[1953] = 24'b000111000001010000000101;
rgb[1954] = 24'b001110000010100100001011;
rgb[1955] = 24'b010101010011111000010001;
rgb[1956] = 24'b011100010101001100010110;
rgb[1957] = 24'b100011010110011100011100;
rgb[1958] = 24'b101010100111110000100010;
rgb[1959] = 24'b110001101001000100100111;
rgb[1960] = 24'b110101111010001000111000;
rgb[1961] = 24'b110111011010111101010100;
rgb[1962] = 24'b111000101011110001110001;
rgb[1963] = 24'b111010001100101010001101;
rgb[1964] = 24'b111011101101011110101010;
rgb[1965] = 24'b111100111110010011000110;
rgb[1966] = 24'b111110011111000111100010;
rgb[1967] = 24'b111111101111111011111111;
rgb[1968] = 24'b000000000000000000000000;
rgb[1969] = 24'b000111010001010100000100;
rgb[1970] = 24'b001110100010101000001001;
rgb[1971] = 24'b010110000011111100001101;
rgb[1972] = 24'b011101010101010000010010;
rgb[1973] = 24'b100100110110100100010110;
rgb[1974] = 24'b101100000111111000011011;
rgb[1975] = 24'b110011101001010000011111;
rgb[1976] = 24'b110111111010010100110000;
rgb[1977] = 24'b111000111011000101001110;
rgb[1978] = 24'b111010001011111001101011;
rgb[1979] = 24'b111011001100101110001001;
rgb[1980] = 24'b111100011101100010100110;
rgb[1981] = 24'b111101011110010111000100;
rgb[1982] = 24'b111110101111001011100001;
rgb[1983] = 24'b111111111111111111111111;
rgb[1984] = 24'b000000000000000000000000;
rgb[1985] = 24'b000111100001010100000011;
rgb[1986] = 24'b001111010010101100000110;
rgb[1987] = 24'b010110110100000000001010;
rgb[1988] = 24'b011110100101011000001101;
rgb[1989] = 24'b100110010110101100010000;
rgb[1990] = 24'b101101111000000100010100;
rgb[1991] = 24'b110101101001011000010111;
rgb[1992] = 24'b111001111010011100101000;
rgb[1993] = 24'b111010101011010001000111;
rgb[1994] = 24'b111011101100000001100101;
rgb[1995] = 24'b111100011100110110000100;
rgb[1996] = 24'b111101001101100110100011;
rgb[1997] = 24'b111110001110011011000001;
rgb[1998] = 24'b111110111111001011100000;
rgb[1999] = 24'b111111111111111111111111;
rgb[2000] = 24'b000000000000000000000000;
rgb[2001] = 24'b000111110001010100000010;
rgb[2002] = 24'b001111110010101100000100;
rgb[2003] = 24'b010111110100000100000110;
rgb[2004] = 24'b011111100101011100001001;
rgb[2005] = 24'b100111100110110100001011;
rgb[2006] = 24'b101111101000001100001101;
rgb[2007] = 24'b110111101001100100001111;
rgb[2008] = 24'b111011111010101000100000;
rgb[2009] = 24'b111100011011011001000000;
rgb[2010] = 24'b111100111100001001100000;
rgb[2011] = 24'b111101011100111010000000;
rgb[2012] = 24'b111110001101101010011111;
rgb[2013] = 24'b111110101110011010111111;
rgb[2014] = 24'b111111001111001011011111;
rgb[2015] = 24'b111111111111111111111111;
rgb[2016] = 24'b000000000000000000000000;
rgb[2017] = 24'b001000000001011000000001;
rgb[2018] = 24'b010000010010110000000010;
rgb[2019] = 24'b011000100100001000000011;
rgb[2020] = 24'b100000110101100100000100;
rgb[2021] = 24'b101001000110111100000101;
rgb[2022] = 24'b110001011000010100000110;
rgb[2023] = 24'b111001101001110000000111;
rgb[2024] = 24'b111101111010110100011000;
rgb[2025] = 24'b111110001011100000111001;
rgb[2026] = 24'b111110011100010001011010;
rgb[2027] = 24'b111110101101000001111011;
rgb[2028] = 24'b111110111101101110011100;
rgb[2029] = 24'b111111001110011110111101;
rgb[2030] = 24'b111111011111001111011110;
rgb[2031] = 24'b111111111111111111111111;
rgb[2032] = 24'b000000000000000000000000;
rgb[2033] = 24'b001000100001011000000000;
rgb[2034] = 24'b010001000010110100000000;
rgb[2035] = 24'b011001100100010000000000;
rgb[2036] = 24'b100010000101101000000000;
rgb[2037] = 24'b101010100111000100000000;
rgb[2038] = 24'b110011001000100000000000;
rgb[2039] = 24'b111011101001111000000000;
rgb[2040] = 24'b111111101010111100010001;
rgb[2041] = 24'b111111111011101100110010;
rgb[2042] = 24'b111111101100011001010101;
rgb[2043] = 24'b111111111101000101110110;
rgb[2044] = 24'b111111111101110110011001;
rgb[2045] = 24'b111111111110100010111011;
rgb[2046] = 24'b111111111111001111011101;
rgb[2047] = 24'b111111111111111111111111;
rgb[2048] = 24'b000000000000000000000000;
rgb[2049] = 24'b000100010001000100010001;
rgb[2050] = 24'b001000100010001000100010;
rgb[2051] = 24'b001100110011001100110011;
rgb[2052] = 24'b010001000100010001000100;
rgb[2053] = 24'b010101010101010101010101;
rgb[2054] = 24'b011001100110011001100110;
rgb[2055] = 24'b011101110111011101110111;
rgb[2056] = 24'b100010001000100010001000;
rgb[2057] = 24'b100110011001100110011001;
rgb[2058] = 24'b101010101010101010101010;
rgb[2059] = 24'b101110111011101110111011;
rgb[2060] = 24'b110011001100110011001100;
rgb[2061] = 24'b110111011101110111011101;
rgb[2062] = 24'b111011101110111011101110;
rgb[2063] = 24'b111111111111111111111111;
rgb[2064] = 24'b000000000000000000000000;
rgb[2065] = 24'b000100100001000100001111;
rgb[2066] = 24'b001001000010001100011111;
rgb[2067] = 24'b001101100011010000101111;
rgb[2068] = 24'b010010000100011000111111;
rgb[2069] = 24'b010110100101011101001111;
rgb[2070] = 24'b011011000110100101011111;
rgb[2071] = 24'b011111100111101101101111;
rgb[2072] = 24'b100011111000110010000000;
rgb[2073] = 24'b100111111001110010010010;
rgb[2074] = 24'b101011111010110010100100;
rgb[2075] = 24'b101111111011110110110110;
rgb[2076] = 24'b110011111100110111001000;
rgb[2077] = 24'b110111111101111011011010;
rgb[2078] = 24'b111011111110111011101100;
rgb[2079] = 24'b111111111111111111111111;
rgb[2080] = 24'b000000000000000000000000;
rgb[2081] = 24'b000100110001001000001110;
rgb[2082] = 24'b001001100010010000011101;
rgb[2083] = 24'b001110010011011000101100;
rgb[2084] = 24'b010011010100100000111010;
rgb[2085] = 24'b011000000101101001001001;
rgb[2086] = 24'b011100110110110101011000;
rgb[2087] = 24'b100001100111111101100111;
rgb[2088] = 24'b100101111001000001111000;
rgb[2089] = 24'b101001101010000010001011;
rgb[2090] = 24'b101101011010111110011110;
rgb[2091] = 24'b110001001011111110110001;
rgb[2092] = 24'b110100101100111111000101;
rgb[2093] = 24'b111000011101111111011000;
rgb[2094] = 24'b111100001110111111101011;
rgb[2095] = 24'b111111111111111111111111;
rgb[2096] = 24'b000000000000000000000000;
rgb[2097] = 24'b000101000001001000001101;
rgb[2098] = 24'b001010000010010100011011;
rgb[2099] = 24'b001111010011100000101000;
rgb[2100] = 24'b010100010100101100110110;
rgb[2101] = 24'b011001010101110101000100;
rgb[2102] = 24'b011110100111000001010001;
rgb[2103] = 24'b100011101000001101011111;
rgb[2104] = 24'b100111111001010001110000;
rgb[2105] = 24'b101011011010001110000100;
rgb[2106] = 24'b101110111011001010011000;
rgb[2107] = 24'b110010001100001010101101;
rgb[2108] = 24'b110101101101000111000001;
rgb[2109] = 24'b111000111110000011010110;
rgb[2110] = 24'b111100011110111111101010;
rgb[2111] = 24'b111111111111111111111111;
rgb[2112] = 24'b000000000000000000000000;
rgb[2113] = 24'b000101010001001100001100;
rgb[2114] = 24'b001010110010011000011000;
rgb[2115] = 24'b010000000011101000100101;
rgb[2116] = 24'b010101100100110100110001;
rgb[2117] = 24'b011010110110000000111110;
rgb[2118] = 24'b100000010111010001001010;
rgb[2119] = 24'b100101101000011101010111;
rgb[2120] = 24'b101001111001100001101000;
rgb[2121] = 24'b101101001010011101111101;
rgb[2122] = 24'b110000001011010110010011;
rgb[2123] = 24'b110011011100010010101000;
rgb[2124] = 24'b110110011101001110111110;
rgb[2125] = 24'b111001101110000111010011;
rgb[2126] = 24'b111100101111000011101001;
rgb[2127] = 24'b111111111111111111111111;
rgb[2128] = 24'b000000000000000000000000;
rgb[2129] = 24'b000101100001001100001011;
rgb[2130] = 24'b001011010010011100010110;
rgb[2131] = 24'b010001000011101100100010;
rgb[2132] = 24'b010110100100111100101101;
rgb[2133] = 24'b011100010110001100111000;
rgb[2134] = 24'b100010000111011101000100;
rgb[2135] = 24'b100111101000101101001111;
rgb[2136] = 24'b101011111001110001100000;
rgb[2137] = 24'b101110111010101001110110;
rgb[2138] = 24'b110001101011100010001101;
rgb[2139] = 24'b110100011100011010100100;
rgb[2140] = 24'b110111011101010010111011;
rgb[2141] = 24'b111010001110001011010001;
rgb[2142] = 24'b111100111111000011101000;
rgb[2143] = 24'b111111111111111111111111;
rgb[2144] = 24'b000000000000000000000000;
rgb[2145] = 24'b000101110001010000001010;
rgb[2146] = 24'b001011110010100100010100;
rgb[2147] = 24'b010001110011110100011110;
rgb[2148] = 24'b010111110101001000101000;
rgb[2149] = 24'b011101100110011000110011;
rgb[2150] = 24'b100011100111101100111101;
rgb[2151] = 24'b101001101000111101000111;
rgb[2152] = 24'b101101111010000001011000;
rgb[2153] = 24'b110000011010111001110000;
rgb[2154] = 24'b110011001011101110000111;
rgb[2155] = 24'b110101101100100110011111;
rgb[2156] = 24'b111000001101011010110111;
rgb[2157] = 24'b111010101110010011001111;
rgb[2158] = 24'b111101001111000111100111;
rgb[2159] = 24'b111111101111111011111111;
rgb[2160] = 24'b000000000000000000000000;
rgb[2161] = 24'b000110000001010100001001;
rgb[2162] = 24'b001100010010101000010010;
rgb[2163] = 24'b010010100011111100011011;
rgb[2164] = 24'b011000110101010000100100;
rgb[2165] = 24'b011111000110100100101101;
rgb[2166] = 24'b100101010111111000110110;
rgb[2167] = 24'b101011101001010000111111;
rgb[2168] = 24'b101111111010010101010000;
rgb[2169] = 24'b110010001011000101101001;
rgb[2170] = 24'b110100011011111010000010;
rgb[2171] = 24'b110110101100101110011011;
rgb[2172] = 24'b111000111101100010110100;
rgb[2173] = 24'b111011001110010111001101;
rgb[2174] = 24'b111101011111001011100110;
rgb[2175] = 24'b111111111111111111111111;
rgb[2176] = 24'b000000000000000000000000;
rgb[2177] = 24'b000110100001010100000111;
rgb[2178] = 24'b001101000010101100001111;
rgb[2179] = 24'b010011100100000100010111;
rgb[2180] = 24'b011010000101011000011111;
rgb[2181] = 24'b100000100110110000100111;
rgb[2182] = 24'b100111001000001000101111;
rgb[2183] = 24'b101101101001100000110111;
rgb[2184] = 24'b110001111010100101001000;
rgb[2185] = 24'b110011111011010101100010;
rgb[2186] = 24'b110101111100000101111100;
rgb[2187] = 24'b110111111100110110010110;
rgb[2188] = 24'b111001111101101010110000;
rgb[2189] = 24'b111011111110011011001010;
rgb[2190] = 24'b111101111111001011100100;
rgb[2191] = 24'b111111101111111011111111;
rgb[2192] = 24'b000000000000000000000000;
rgb[2193] = 24'b000110110001011000000110;
rgb[2194] = 24'b001101100010110000001101;
rgb[2195] = 24'b010100010100001100010100;
rgb[2196] = 24'b011011000101100100011011;
rgb[2197] = 24'b100010000110111100100001;
rgb[2198] = 24'b101000111000011000101000;
rgb[2199] = 24'b101111101001110000101111;
rgb[2200] = 24'b110011111010110101000000;
rgb[2201] = 24'b110101101011100101011011;
rgb[2202] = 24'b110111011100010001110110;
rgb[2203] = 24'b111000111101000010010010;
rgb[2204] = 24'b111010101101110010101101;
rgb[2205] = 24'b111100011110011111001000;
rgb[2206] = 24'b111110001111001111100011;
rgb[2207] = 24'b111111111111111111111111;
rgb[2208] = 24'b000000000000000000000000;
rgb[2209] = 24'b000111000001011000000101;
rgb[2210] = 24'b001110000010110100001011;
rgb[2211] = 24'b010101010100010000010001;
rgb[2212] = 24'b011100010101101100010110;
rgb[2213] = 24'b100011010111001000011100;
rgb[2214] = 24'b101010101000100100100010;
rgb[2215] = 24'b110001101010000000100111;
rgb[2216] = 24'b110101111011000100111000;
rgb[2217] = 24'b110111011011110001010100;
rgb[2218] = 24'b111000101100011101110001;
rgb[2219] = 24'b111010001101001010001101;
rgb[2220] = 24'b111011101101110110101010;
rgb[2221] = 24'b111100111110100011000110;
rgb[2222] = 24'b111110011111001111100010;
rgb[2223] = 24'b111111101111111011111111;
rgb[2224] = 24'b000000000000000000000000;
rgb[2225] = 24'b000111010001011100000100;
rgb[2226] = 24'b001110100010111100001001;
rgb[2227] = 24'b010110000100011000001101;
rgb[2228] = 24'b011101010101111000010010;
rgb[2229] = 24'b100100110111010100010110;
rgb[2230] = 24'b101100001000110100011011;
rgb[2231] = 24'b110011101010010000011111;
rgb[2232] = 24'b110111111011010100110000;
rgb[2233] = 24'b111000111100000001001110;
rgb[2234] = 24'b111010001100101001101011;
rgb[2235] = 24'b111011001101010110001001;
rgb[2236] = 24'b111100011101111110100110;
rgb[2237] = 24'b111101011110101011000100;
rgb[2238] = 24'b111110101111010011100001;
rgb[2239] = 24'b111111111111111111111111;
rgb[2240] = 24'b000000000000000000000000;
rgb[2241] = 24'b000111100001100000000011;
rgb[2242] = 24'b001111010011000000000110;
rgb[2243] = 24'b010110110100100000001010;
rgb[2244] = 24'b011110100110000000001101;
rgb[2245] = 24'b100110010111100000010000;
rgb[2246] = 24'b101101111001000000010100;
rgb[2247] = 24'b110101101010100000010111;
rgb[2248] = 24'b111001111011100100101000;
rgb[2249] = 24'b111010101100001101000111;
rgb[2250] = 24'b111011101100110101100101;
rgb[2251] = 24'b111100011101011110000100;
rgb[2252] = 24'b111101001110000110100011;
rgb[2253] = 24'b111110001110101111000001;
rgb[2254] = 24'b111110111111010111100000;
rgb[2255] = 24'b111111111111111111111111;
rgb[2256] = 24'b000000000000000000000000;
rgb[2257] = 24'b000111110001100000000010;
rgb[2258] = 24'b001111110011000100000100;
rgb[2259] = 24'b010111110100101000000110;
rgb[2260] = 24'b011111100110001000001001;
rgb[2261] = 24'b100111100111101100001011;
rgb[2262] = 24'b101111101001010000001101;
rgb[2263] = 24'b110111101010110100001111;
rgb[2264] = 24'b111011111011111000100000;
rgb[2265] = 24'b111100011100011101000000;
rgb[2266] = 24'b111100111101000001100000;
rgb[2267] = 24'b111101011101100110000000;
rgb[2268] = 24'b111110001110001110011111;
rgb[2269] = 24'b111110101110110010111111;
rgb[2270] = 24'b111111001111010111011111;
rgb[2271] = 24'b111111111111111111111111;
rgb[2272] = 24'b000000000000000000000000;
rgb[2273] = 24'b001000000001100100000001;
rgb[2274] = 24'b010000010011001000000010;
rgb[2275] = 24'b011000100100101100000011;
rgb[2276] = 24'b100000110110010100000100;
rgb[2277] = 24'b101001000111111000000101;
rgb[2278] = 24'b110001011001011100000110;
rgb[2279] = 24'b111001101011000100000111;
rgb[2280] = 24'b111101111100001000011000;
rgb[2281] = 24'b111110001100101000111001;
rgb[2282] = 24'b111110011101001101011010;
rgb[2283] = 24'b111110101101110001111011;
rgb[2284] = 24'b111110111110010010011100;
rgb[2285] = 24'b111111001110110110111101;
rgb[2286] = 24'b111111011111011011011110;
rgb[2287] = 24'b111111111111111111111111;
rgb[2288] = 24'b000000000000000000000000;
rgb[2289] = 24'b001000100001100100000000;
rgb[2290] = 24'b010001000011001100000000;
rgb[2291] = 24'b011001100100110100000000;
rgb[2292] = 24'b100010000110011100000000;
rgb[2293] = 24'b101010101000000100000000;
rgb[2294] = 24'b110011001001101100000000;
rgb[2295] = 24'b111011101011010100000000;
rgb[2296] = 24'b111111101100011000010001;
rgb[2297] = 24'b111111111100111000110010;
rgb[2298] = 24'b111111101101011001010101;
rgb[2299] = 24'b111111111101111001110110;
rgb[2300] = 24'b111111111110011010011001;
rgb[2301] = 24'b111111111110111010111011;
rgb[2302] = 24'b111111111111011011011101;
rgb[2303] = 24'b111111111111111111111111;
rgb[2304] = 24'b000000000000000000000000;
rgb[2305] = 24'b000100010001000100010001;
rgb[2306] = 24'b001000100010001000100010;
rgb[2307] = 24'b001100110011001100110011;
rgb[2308] = 24'b010001000100010001000100;
rgb[2309] = 24'b010101010101010101010101;
rgb[2310] = 24'b011001100110011001100110;
rgb[2311] = 24'b011101110111011101110111;
rgb[2312] = 24'b100010001000100010001000;
rgb[2313] = 24'b100110011001100110011001;
rgb[2314] = 24'b101010101010101010101010;
rgb[2315] = 24'b101110111011101110111011;
rgb[2316] = 24'b110011001100110011001100;
rgb[2317] = 24'b110111011101110111011101;
rgb[2318] = 24'b111011101110111011101110;
rgb[2319] = 24'b111111111111111111111111;
rgb[2320] = 24'b000000000000000000000000;
rgb[2321] = 24'b000100100001000100001111;
rgb[2322] = 24'b001001000010001100011111;
rgb[2323] = 24'b001101100011010100101111;
rgb[2324] = 24'b010010000100011100111111;
rgb[2325] = 24'b010110100101100101001111;
rgb[2326] = 24'b011011000110101001011111;
rgb[2327] = 24'b011111100111110001101111;
rgb[2328] = 24'b100011111000110110000000;
rgb[2329] = 24'b100111111001110110010010;
rgb[2330] = 24'b101011111010111010100100;
rgb[2331] = 24'b101111111011111010110110;
rgb[2332] = 24'b110011111100111011001000;
rgb[2333] = 24'b110111111101111011011010;
rgb[2334] = 24'b111011111110111011101100;
rgb[2335] = 24'b111111111111111111111111;
rgb[2336] = 24'b000000000000000000000000;
rgb[2337] = 24'b000100110001001000001110;
rgb[2338] = 24'b001001100010010100011101;
rgb[2339] = 24'b001110010011011100101100;
rgb[2340] = 24'b010011010100101000111010;
rgb[2341] = 24'b011000000101110101001001;
rgb[2342] = 24'b011100110110111101011000;
rgb[2343] = 24'b100001101000001001100111;
rgb[2344] = 24'b100101111001001101111000;
rgb[2345] = 24'b101001101010001010001011;
rgb[2346] = 24'b101101011011001010011110;
rgb[2347] = 24'b110001001100000110110001;
rgb[2348] = 24'b110100101101000011000101;
rgb[2349] = 24'b111000011110000011011000;
rgb[2350] = 24'b111100001110111111101011;
rgb[2351] = 24'b111111111111111111111111;
rgb[2352] = 24'b000000000000000000000000;
rgb[2353] = 24'b000101000001001100001101;
rgb[2354] = 24'b001010000010011000011011;
rgb[2355] = 24'b001111010011101000101000;
rgb[2356] = 24'b010100010100110100110110;
rgb[2357] = 24'b011001010110000101000100;
rgb[2358] = 24'b011110100111010001010001;
rgb[2359] = 24'b100011101000100001011111;
rgb[2360] = 24'b100111111001100101110000;
rgb[2361] = 24'b101011011010011110000100;
rgb[2362] = 24'b101110111011011010011000;
rgb[2363] = 24'b110010001100010010101101;
rgb[2364] = 24'b110101101101001111000001;
rgb[2365] = 24'b111000111110000111010110;
rgb[2366] = 24'b111100011111000011101010;
rgb[2367] = 24'b111111111111111111111111;
rgb[2368] = 24'b000000000000000000000000;
rgb[2369] = 24'b000101010001010000001100;
rgb[2370] = 24'b001010110010100000011000;
rgb[2371] = 24'b010000000011110000100101;
rgb[2372] = 24'b010101100101000000110001;
rgb[2373] = 24'b011010110110010100111110;
rgb[2374] = 24'b100000010111100101001010;
rgb[2375] = 24'b100101101000110101010111;
rgb[2376] = 24'b101001111001111001101000;
rgb[2377] = 24'b101101001010110001111101;
rgb[2378] = 24'b110000001011101010010011;
rgb[2379] = 24'b110011011100011110101000;
rgb[2380] = 24'b110110011101010110111110;
rgb[2381] = 24'b111001101110001111010011;
rgb[2382] = 24'b111100101111000111101001;
rgb[2383] = 24'b111111111111111111111111;
rgb[2384] = 24'b000000000000000000000000;
rgb[2385] = 24'b000101100001010100001011;
rgb[2386] = 24'b001011010010101000010110;
rgb[2387] = 24'b010001000011111100100010;
rgb[2388] = 24'b010110100101010000101101;
rgb[2389] = 24'b011100010110100100111000;
rgb[2390] = 24'b100010000111111001000100;
rgb[2391] = 24'b100111101001001101001111;
rgb[2392] = 24'b101011111010010001100000;
rgb[2393] = 24'b101110111011000101110110;
rgb[2394] = 24'b110001101011111010001101;
rgb[2395] = 24'b110100011100101110100100;
rgb[2396] = 24'b110111011101100010111011;
rgb[2397] = 24'b111010001110010111010001;
rgb[2398] = 24'b111100111111001011101000;
rgb[2399] = 24'b111111111111111111111111;
rgb[2400] = 24'b000000000000000000000000;
rgb[2401] = 24'b000101110001010100001010;
rgb[2402] = 24'b001011110010101100010100;
rgb[2403] = 24'b010001110100000100011110;
rgb[2404] = 24'b010111110101011100101000;
rgb[2405] = 24'b011101100110110100110011;
rgb[2406] = 24'b100011101000001100111101;
rgb[2407] = 24'b101001101001100101000111;
rgb[2408] = 24'b101101111010101001011000;
rgb[2409] = 24'b110000011011011001110000;
rgb[2410] = 24'b110011001100001010000111;
rgb[2411] = 24'b110101101100111010011111;
rgb[2412] = 24'b111000001101101010110111;
rgb[2413] = 24'b111010101110011011001111;
rgb[2414] = 24'b111101001111001011100111;
rgb[2415] = 24'b111111101111111011111111;
rgb[2416] = 24'b000000000000000000000000;
rgb[2417] = 24'b000110000001011000001001;
rgb[2418] = 24'b001100010010110100010010;
rgb[2419] = 24'b010010100100010000011011;
rgb[2420] = 24'b011000110101101000100100;
rgb[2421] = 24'b011111000111000100101101;
rgb[2422] = 24'b100101011000100000110110;
rgb[2423] = 24'b101011101001111000111111;
rgb[2424] = 24'b101111111010111101010000;
rgb[2425] = 24'b110010001011101101101001;
rgb[2426] = 24'b110100011100011010000010;
rgb[2427] = 24'b110110101101000110011011;
rgb[2428] = 24'b111000111101110110110100;
rgb[2429] = 24'b111011001110100011001101;
rgb[2430] = 24'b111101011111001111100110;
rgb[2431] = 24'b111111111111111111111111;
rgb[2432] = 24'b000000000000000000000000;
rgb[2433] = 24'b000110100001011100000111;
rgb[2434] = 24'b001101000010111000001111;
rgb[2435] = 24'b010011100100011000010111;
rgb[2436] = 24'b011010000101110100011111;
rgb[2437] = 24'b100000100111010100100111;
rgb[2438] = 24'b100111001000110000101111;
rgb[2439] = 24'b101101101010010000110111;
rgb[2440] = 24'b110001111011010101001000;
rgb[2441] = 24'b110011111011111101100010;
rgb[2442] = 24'b110101111100101001111100;
rgb[2443] = 24'b110111111101010010010110;
rgb[2444] = 24'b111001111101111110110000;
rgb[2445] = 24'b111011111110100111001010;
rgb[2446] = 24'b111101111111010011100100;
rgb[2447] = 24'b111111101111111011111111;
rgb[2448] = 24'b000000000000000000000000;
rgb[2449] = 24'b000110110001100000000110;
rgb[2450] = 24'b001101100011000000001101;
rgb[2451] = 24'b010100010100100000010100;
rgb[2452] = 24'b011011000110000100011011;
rgb[2453] = 24'b100010000111100100100001;
rgb[2454] = 24'b101000111001000100101000;
rgb[2455] = 24'b101111101010101000101111;
rgb[2456] = 24'b110011111011101101000000;
rgb[2457] = 24'b110101101100010001011011;
rgb[2458] = 24'b110111011100111001110110;
rgb[2459] = 24'b111000111101100010010010;
rgb[2460] = 24'b111010101110000110101101;
rgb[2461] = 24'b111100011110101111001000;
rgb[2462] = 24'b111110001111010111100011;
rgb[2463] = 24'b111111111111111111111111;
rgb[2464] = 24'b000000000000000000000000;
rgb[2465] = 24'b000111000001100100000101;
rgb[2466] = 24'b001110000011001000001011;
rgb[2467] = 24'b010101010100101100010001;
rgb[2468] = 24'b011100010110010000010110;
rgb[2469] = 24'b100011010111110100011100;
rgb[2470] = 24'b101010101001011000100010;
rgb[2471] = 24'b110001101010111100100111;
rgb[2472] = 24'b110101111100000000111000;
rgb[2473] = 24'b110111011100100101010100;
rgb[2474] = 24'b111000101101001001110001;
rgb[2475] = 24'b111010001101101110001101;
rgb[2476] = 24'b111011101110010010101010;
rgb[2477] = 24'b111100111110110111000110;
rgb[2478] = 24'b111110011111011011100010;
rgb[2479] = 24'b111111101111111011111111;
rgb[2480] = 24'b000000000000000000000000;
rgb[2481] = 24'b000111010001100100000100;
rgb[2482] = 24'b001110100011001100001001;
rgb[2483] = 24'b010110000100110100001101;
rgb[2484] = 24'b011101010110011100010010;
rgb[2485] = 24'b100100111000000100010110;
rgb[2486] = 24'b101100001001101100011011;
rgb[2487] = 24'b110011101011010100011111;
rgb[2488] = 24'b110111111100011000110000;
rgb[2489] = 24'b111000111100111001001110;
rgb[2490] = 24'b111010001101011001101011;
rgb[2491] = 24'b111011001101111010001001;
rgb[2492] = 24'b111100011110011010100110;
rgb[2493] = 24'b111101011110111011000100;
rgb[2494] = 24'b111110101111011011100001;
rgb[2495] = 24'b111111111111111111111111;
rgb[2496] = 24'b000000000000000000000000;
rgb[2497] = 24'b000111100001101000000011;
rgb[2498] = 24'b001111010011010100000110;
rgb[2499] = 24'b010110110101000000001010;
rgb[2500] = 24'b011110100110101000001101;
rgb[2501] = 24'b100110011000010100010000;
rgb[2502] = 24'b101101111010000000010100;
rgb[2503] = 24'b110101101011101100010111;
rgb[2504] = 24'b111001111100110000101000;
rgb[2505] = 24'b111010101101001101000111;
rgb[2506] = 24'b111011101101101001100101;
rgb[2507] = 24'b111100011110000110000100;
rgb[2508] = 24'b111101001110100110100011;
rgb[2509] = 24'b111110001111000011000001;
rgb[2510] = 24'b111110111111011111100000;
rgb[2511] = 24'b111111111111111111111111;
rgb[2512] = 24'b000000000000000000000000;
rgb[2513] = 24'b000111110001101100000010;
rgb[2514] = 24'b001111110011011100000100;
rgb[2515] = 24'b010111110101001000000110;
rgb[2516] = 24'b011111100110111000001001;
rgb[2517] = 24'b100111101000100100001011;
rgb[2518] = 24'b101111101010010100001101;
rgb[2519] = 24'b110111101100000000001111;
rgb[2520] = 24'b111011111101000100100000;
rgb[2521] = 24'b111100011101100001000000;
rgb[2522] = 24'b111100111101111001100000;
rgb[2523] = 24'b111101011110010110000000;
rgb[2524] = 24'b111110001110101110011111;
rgb[2525] = 24'b111110101111001010111111;
rgb[2526] = 24'b111111001111100011011111;
rgb[2527] = 24'b111111111111111111111111;
rgb[2528] = 24'b000000000000000000000000;
rgb[2529] = 24'b001000000001110000000001;
rgb[2530] = 24'b010000010011100000000010;
rgb[2531] = 24'b011000100101010100000011;
rgb[2532] = 24'b100000110111000100000100;
rgb[2533] = 24'b101001001000110100000101;
rgb[2534] = 24'b110001011010101000000110;
rgb[2535] = 24'b111001101100011000000111;
rgb[2536] = 24'b111101111101011100011000;
rgb[2537] = 24'b111110001101110000111001;
rgb[2538] = 24'b111110011110001001011010;
rgb[2539] = 24'b111110101110100001111011;
rgb[2540] = 24'b111110111110111010011100;
rgb[2541] = 24'b111111001111001110111101;
rgb[2542] = 24'b111111011111100111011110;
rgb[2543] = 24'b111111111111111111111111;
rgb[2544] = 24'b000000000000000000000000;
rgb[2545] = 24'b001000100001110100000000;
rgb[2546] = 24'b010001000011101000000000;
rgb[2547] = 24'b011001100101011100000000;
rgb[2548] = 24'b100010000111010000000000;
rgb[2549] = 24'b101010101001000100000000;
rgb[2550] = 24'b110011001010111000000000;
rgb[2551] = 24'b111011101100110000000000;
rgb[2552] = 24'b111111101101110000010001;
rgb[2553] = 24'b111111111110000100110010;
rgb[2554] = 24'b111111101110011001010101;
rgb[2555] = 24'b111111111110101101110110;
rgb[2556] = 24'b111111111111000010011001;
rgb[2557] = 24'b111111111111010110111011;
rgb[2558] = 24'b111111111111101011011101;
rgb[2559] = 24'b111111111111111111111111;
rgb[2560] = 24'b000000000000000000000000;
rgb[2561] = 24'b000100010001000100010001;
rgb[2562] = 24'b001000100010001000100010;
rgb[2563] = 24'b001100110011001100110011;
rgb[2564] = 24'b010001000100010001000100;
rgb[2565] = 24'b010101010101010101010101;
rgb[2566] = 24'b011001100110011001100110;
rgb[2567] = 24'b011101110111011101110111;
rgb[2568] = 24'b100010001000100010001000;
rgb[2569] = 24'b100110011001100110011001;
rgb[2570] = 24'b101010101010101010101010;
rgb[2571] = 24'b101110111011101110111011;
rgb[2572] = 24'b110011001100110011001100;
rgb[2573] = 24'b110111011101110111011101;
rgb[2574] = 24'b111011101110111011101110;
rgb[2575] = 24'b111111111111111111111111;
rgb[2576] = 24'b000000000000000000000000;
rgb[2577] = 24'b000100100001001000001111;
rgb[2578] = 24'b001001000010010000011111;
rgb[2579] = 24'b001101100011011000101111;
rgb[2580] = 24'b010010000100100000111111;
rgb[2581] = 24'b010110100101101001001111;
rgb[2582] = 24'b011011000110110001011111;
rgb[2583] = 24'b011111100111111001101111;
rgb[2584] = 24'b100011111000111110000000;
rgb[2585] = 24'b100111111001111110010010;
rgb[2586] = 24'b101011111010111110100100;
rgb[2587] = 24'b101111111011111110110110;
rgb[2588] = 24'b110011111100111111001000;
rgb[2589] = 24'b110111111101111111011010;
rgb[2590] = 24'b111011111110111111101100;
rgb[2591] = 24'b111111111111111111111111;
rgb[2592] = 24'b000000000000000000000000;
rgb[2593] = 24'b000100110001001100001110;
rgb[2594] = 24'b001001100010011000011101;
rgb[2595] = 24'b001110010011100100101100;
rgb[2596] = 24'b010011010100110000111010;
rgb[2597] = 24'b011000000101111101001001;
rgb[2598] = 24'b011100110111001001011000;
rgb[2599] = 24'b100001101000010101100111;
rgb[2600] = 24'b100101111001011001111000;
rgb[2601] = 24'b101001101010010110001011;
rgb[2602] = 24'b101101011011010010011110;
rgb[2603] = 24'b110001001100001110110001;
rgb[2604] = 24'b110100101101001011000101;
rgb[2605] = 24'b111000011110000111011000;
rgb[2606] = 24'b111100001111000011101011;
rgb[2607] = 24'b111111111111111111111111;
rgb[2608] = 24'b000000000000000000000000;
rgb[2609] = 24'b000101000001010000001101;
rgb[2610] = 24'b001010000010100000011011;
rgb[2611] = 24'b001111010011110000101000;
rgb[2612] = 24'b010100010101000000110110;
rgb[2613] = 24'b011001010110010001000100;
rgb[2614] = 24'b011110100111100001010001;
rgb[2615] = 24'b100011101000110001011111;
rgb[2616] = 24'b100111111001110101110000;
rgb[2617] = 24'b101011011010101110000100;
rgb[2618] = 24'b101110111011100110011000;
rgb[2619] = 24'b110010001100011110101101;
rgb[2620] = 24'b110101101101010111000001;
rgb[2621] = 24'b111000111110001111010110;
rgb[2622] = 24'b111100011111000111101010;
rgb[2623] = 24'b111111111111111111111111;
rgb[2624] = 24'b000000000000000000000000;
rgb[2625] = 24'b000101010001010100001100;
rgb[2626] = 24'b001010110010101000011000;
rgb[2627] = 24'b010000000011111100100101;
rgb[2628] = 24'b010101100101010000110001;
rgb[2629] = 24'b011010110110100100111110;
rgb[2630] = 24'b100000010111111001001010;
rgb[2631] = 24'b100101101001001101010111;
rgb[2632] = 24'b101001111010010001101000;
rgb[2633] = 24'b101101001011000101111101;
rgb[2634] = 24'b110000001011111010010011;
rgb[2635] = 24'b110011011100101110101000;
rgb[2636] = 24'b110110011101100010111110;
rgb[2637] = 24'b111001101110010111010011;
rgb[2638] = 24'b111100101111001011101001;
rgb[2639] = 24'b111111111111111111111111;
rgb[2640] = 24'b000000000000000000000000;
rgb[2641] = 24'b000101100001011000001011;
rgb[2642] = 24'b001011010010110000010110;
rgb[2643] = 24'b010001000100001000100010;
rgb[2644] = 24'b010110100101100000101101;
rgb[2645] = 24'b011100010110111000111000;
rgb[2646] = 24'b100010001000010001000100;
rgb[2647] = 24'b100111101001101001001111;
rgb[2648] = 24'b101011111010101101100000;
rgb[2649] = 24'b101110111011011101110110;
rgb[2650] = 24'b110001101100001110001101;
rgb[2651] = 24'b110100011100111110100100;
rgb[2652] = 24'b110111011101101110111011;
rgb[2653] = 24'b111010001110011111010001;
rgb[2654] = 24'b111100111111001111101000;
rgb[2655] = 24'b111111111111111111111111;
rgb[2656] = 24'b000000000000000000000000;
rgb[2657] = 24'b000101110001011100001010;
rgb[2658] = 24'b001011110010111000010100;
rgb[2659] = 24'b010001110100010100011110;
rgb[2660] = 24'b010111110101110000101000;
rgb[2661] = 24'b011101100111001100110011;
rgb[2662] = 24'b100011101000101000111101;
rgb[2663] = 24'b101001101010001001000111;
rgb[2664] = 24'b101101111011001101011000;
rgb[2665] = 24'b110000011011110101110000;
rgb[2666] = 24'b110011001100100010000111;
rgb[2667] = 24'b110101101101001110011111;
rgb[2668] = 24'b111000001101111010110111;
rgb[2669] = 24'b111010101110100111001111;
rgb[2670] = 24'b111101001111010011100111;
rgb[2671] = 24'b111111101111111011111111;
rgb[2672] = 24'b000000000000000000000000;
rgb[2673] = 24'b000110000001100000001001;
rgb[2674] = 24'b001100010011000000010010;
rgb[2675] = 24'b010010100100100000011011;
rgb[2676] = 24'b011000110110000000100100;
rgb[2677] = 24'b011111000111100000101101;
rgb[2678] = 24'b100101011001000100110110;
rgb[2679] = 24'b101011101010100100111111;
rgb[2680] = 24'b101111111011101001010000;
rgb[2681] = 24'b110010001100010001101001;
rgb[2682] = 24'b110100011100110110000010;
rgb[2683] = 24'b110110101101011110011011;
rgb[2684] = 24'b111000111110000110110100;
rgb[2685] = 24'b111011001110101111001101;
rgb[2686] = 24'b111101011111010111100110;
rgb[2687] = 24'b111111111111111111111111;
rgb[2688] = 24'b000000000000000000000000;
rgb[2689] = 24'b000110100001100100000111;
rgb[2690] = 24'b001101000011001000001111;
rgb[2691] = 24'b010011100100101100010111;
rgb[2692] = 24'b011010000110010000011111;
rgb[2693] = 24'b100000100111111000100111;
rgb[2694] = 24'b100111001001011100101111;
rgb[2695] = 24'b101101101011000000110111;
rgb[2696] = 24'b110001111100000101001000;
rgb[2697] = 24'b110011111100101001100010;
rgb[2698] = 24'b110101111101001101111100;
rgb[2699] = 24'b110111111101101110010110;
rgb[2700] = 24'b111001111110010010110000;
rgb[2701] = 24'b111011111110110111001010;
rgb[2702] = 24'b111101111111011011100100;
rgb[2703] = 24'b111111101111111011111111;
rgb[2704] = 24'b000000000000000000000000;
rgb[2705] = 24'b000110110001101000000110;
rgb[2706] = 24'b001101100011010000001101;
rgb[2707] = 24'b010100010100111000010100;
rgb[2708] = 24'b011011000110100000011011;
rgb[2709] = 24'b100010001000001100100001;
rgb[2710] = 24'b101000111001110100101000;
rgb[2711] = 24'b101111101011011100101111;
rgb[2712] = 24'b110011111100100001000000;
rgb[2713] = 24'b110101101101000001011011;
rgb[2714] = 24'b110111011101100001110110;
rgb[2715] = 24'b111000111101111110010010;
rgb[2716] = 24'b111010101110011110101101;
rgb[2717] = 24'b111100011110111111001000;
rgb[2718] = 24'b111110001111011111100011;
rgb[2719] = 24'b111111111111111111111111;
rgb[2720] = 24'b000000000000000000000000;
rgb[2721] = 24'b000111000001101100000101;
rgb[2722] = 24'b001110000011011000001011;
rgb[2723] = 24'b010101010101000100010001;
rgb[2724] = 24'b011100010110110100010110;
rgb[2725] = 24'b100011011000100000011100;
rgb[2726] = 24'b101010101010001100100010;
rgb[2727] = 24'b110001101011111000100111;
rgb[2728] = 24'b110101111100111100111000;
rgb[2729] = 24'b110111011101011001010100;
rgb[2730] = 24'b111000101101110101110001;
rgb[2731] = 24'b111010001110010010001101;
rgb[2732] = 24'b111011101110101010101010;
rgb[2733] = 24'b111100111111000111000110;
rgb[2734] = 24'b111110011111100011100010;
rgb[2735] = 24'b111111101111111011111111;
rgb[2736] = 24'b000000000000000000000000;
rgb[2737] = 24'b000111010001110000000100;
rgb[2738] = 24'b001110100011100000001001;
rgb[2739] = 24'b010110000101010000001101;
rgb[2740] = 24'b011101010111000100010010;
rgb[2741] = 24'b100100111000110100010110;
rgb[2742] = 24'b101100001010100100011011;
rgb[2743] = 24'b110011101100010100011111;
rgb[2744] = 24'b110111111101011000110000;
rgb[2745] = 24'b111000111101110001001110;
rgb[2746] = 24'b111010001110001001101011;
rgb[2747] = 24'b111011001110100010001001;
rgb[2748] = 24'b111100011110110110100110;
rgb[2749] = 24'b111101011111001111000100;
rgb[2750] = 24'b111110101111100111100001;
rgb[2751] = 24'b111111111111111111111111;
rgb[2752] = 24'b000000000000000000000000;
rgb[2753] = 24'b000111100001110100000011;
rgb[2754] = 24'b001111010011101000000110;
rgb[2755] = 24'b010110110101011100001010;
rgb[2756] = 24'b011110100111010100001101;
rgb[2757] = 24'b100110011001001000010000;
rgb[2758] = 24'b101101111010111100010100;
rgb[2759] = 24'b110101101100110100010111;
rgb[2760] = 24'b111001111101111000101000;
rgb[2761] = 24'b111010101110001001000111;
rgb[2762] = 24'b111011101110011101100101;
rgb[2763] = 24'b111100011110110010000100;
rgb[2764] = 24'b111101001111000010100011;
rgb[2765] = 24'b111110001111010111000001;
rgb[2766] = 24'b111110111111101011100000;
rgb[2767] = 24'b111111111111111111111111;
rgb[2768] = 24'b000000000000000000000000;
rgb[2769] = 24'b000111110001111000000010;
rgb[2770] = 24'b001111110011110000000100;
rgb[2771] = 24'b010111110101101000000110;
rgb[2772] = 24'b011111100111100100001001;
rgb[2773] = 24'b100111101001011100001011;
rgb[2774] = 24'b101111101011010100001101;
rgb[2775] = 24'b110111101101010000001111;
rgb[2776] = 24'b111011111110010100100000;
rgb[2777] = 24'b111100011110100001000000;
rgb[2778] = 24'b111100111110110001100000;
rgb[2779] = 24'b111101011111000010000000;
rgb[2780] = 24'b111110001111001110011111;
rgb[2781] = 24'b111110101111011110111111;
rgb[2782] = 24'b111111001111101111011111;
rgb[2783] = 24'b111111111111111111111111;
rgb[2784] = 24'b000000000000000000000000;
rgb[2785] = 24'b001000000001111100000001;
rgb[2786] = 24'b010000010011111000000010;
rgb[2787] = 24'b011000100101111000000011;
rgb[2788] = 24'b100000110111110100000100;
rgb[2789] = 24'b101001001001110000000101;
rgb[2790] = 24'b110001011011110000000110;
rgb[2791] = 24'b111001101101101100000111;
rgb[2792] = 24'b111101111110110000011000;
rgb[2793] = 24'b111110001110111100111001;
rgb[2794] = 24'b111110011111000101011010;
rgb[2795] = 24'b111110101111010001111011;
rgb[2796] = 24'b111110111111011110011100;
rgb[2797] = 24'b111111001111100110111101;
rgb[2798] = 24'b111111011111110011011110;
rgb[2799] = 24'b111111111111111111111111;
rgb[2800] = 24'b000000000000000000000000;
rgb[2801] = 24'b001000100010000000000000;
rgb[2802] = 24'b010001000100000000000000;
rgb[2803] = 24'b011001100110000100000000;
rgb[2804] = 24'b100010001000000100000000;
rgb[2805] = 24'b101010101010000100000000;
rgb[2806] = 24'b110011001100001000000000;
rgb[2807] = 24'b111011101110001000000000;
rgb[2808] = 24'b111111101111001100010001;
rgb[2809] = 24'b111111111111010100110010;
rgb[2810] = 24'b111111101111011001010101;
rgb[2811] = 24'b111111111111100001110110;
rgb[2812] = 24'b111111111111101010011001;
rgb[2813] = 24'b111111111111101110111011;
rgb[2814] = 24'b111111111111110111011101;
rgb[2815] = 24'b111111111111111111111111;
rgb[2816] = 24'b000000000000000000000000;
rgb[2817] = 24'b000100010001000100010001;
rgb[2818] = 24'b001000100010001000100010;
rgb[2819] = 24'b001100110011001100110011;
rgb[2820] = 24'b010001000100010001000100;
rgb[2821] = 24'b010101010101010101010101;
rgb[2822] = 24'b011001100110011001100110;
rgb[2823] = 24'b011101110111011101110111;
rgb[2824] = 24'b100010001000100010001000;
rgb[2825] = 24'b100110011001100110011001;
rgb[2826] = 24'b101010101010101010101010;
rgb[2827] = 24'b101110111011101110111011;
rgb[2828] = 24'b110011001100110011001100;
rgb[2829] = 24'b110111011101110111011101;
rgb[2830] = 24'b111011101110111011101110;
rgb[2831] = 24'b111111111111111111111111;
rgb[2832] = 24'b000000000000000000000000;
rgb[2833] = 24'b000100100001001000001111;
rgb[2834] = 24'b001001000010010000011111;
rgb[2835] = 24'b001101100011011000101111;
rgb[2836] = 24'b010010000100100000111111;
rgb[2837] = 24'b010110100101101001001111;
rgb[2838] = 24'b011011000110110001011111;
rgb[2839] = 24'b011111100111111001101111;
rgb[2840] = 24'b100011111000111110000000;
rgb[2841] = 24'b100111111001111110010010;
rgb[2842] = 24'b101011111010111110100100;
rgb[2843] = 24'b101111111011111110110110;
rgb[2844] = 24'b110011111100111111001000;
rgb[2845] = 24'b110111111101111111011010;
rgb[2846] = 24'b111011111110111111101100;
rgb[2847] = 24'b111111111111111111111111;
rgb[2848] = 24'b000000000000000000000000;
rgb[2849] = 24'b000100110001001100001110;
rgb[2850] = 24'b001001100010011000011101;
rgb[2851] = 24'b001110010011100100101100;
rgb[2852] = 24'b010011000100110100111010;
rgb[2853] = 24'b010111110110000001001001;
rgb[2854] = 24'b011100100111001101011000;
rgb[2855] = 24'b100001011000011001100111;
rgb[2856] = 24'b100101101001011101111000;
rgb[2857] = 24'b101001011010011010001011;
rgb[2858] = 24'b101101001011010110011110;
rgb[2859] = 24'b110000111100010010110001;
rgb[2860] = 24'b110100101101001011000101;
rgb[2861] = 24'b111000011110000111011000;
rgb[2862] = 24'b111100001111000011101011;
rgb[2863] = 24'b111111111111111111111111;
rgb[2864] = 24'b000000000000000000000000;
rgb[2865] = 24'b000101000001010000001101;
rgb[2866] = 24'b001010000010100000011011;
rgb[2867] = 24'b001111000011110100101000;
rgb[2868] = 24'b010100000101000100110110;
rgb[2869] = 24'b011001000110010101000100;
rgb[2870] = 24'b011110000111101001010001;
rgb[2871] = 24'b100011001000111001011111;
rgb[2872] = 24'b100111011001111101110000;
rgb[2873] = 24'b101010111010110110000100;
rgb[2874] = 24'b101110011011101110011000;
rgb[2875] = 24'b110001111100100010101101;
rgb[2876] = 24'b110101011101011011000001;
rgb[2877] = 24'b111000111110001111010110;
rgb[2878] = 24'b111100011111000111101010;
rgb[2879] = 24'b111111111111111111111111;
rgb[2880] = 24'b000000000000000000000000;
rgb[2881] = 24'b000101010001010100001100;
rgb[2882] = 24'b001010100010101100011000;
rgb[2883] = 24'b001111110100000000100101;
rgb[2884] = 24'b010101000101011000110001;
rgb[2885] = 24'b011010010110101100111110;
rgb[2886] = 24'b011111101000000101001010;
rgb[2887] = 24'b100100111001011001010111;
rgb[2888] = 24'b101001001010011101101000;
rgb[2889] = 24'b101100011011010001111101;
rgb[2890] = 24'b101111101100000010010011;
rgb[2891] = 24'b110010111100110110101000;
rgb[2892] = 24'b110110001101100110111110;
rgb[2893] = 24'b111001011110011011010011;
rgb[2894] = 24'b111100101111001011101001;
rgb[2895] = 24'b111111111111111111111111;
rgb[2896] = 24'b000000000000000000000000;
rgb[2897] = 24'b000101100001011000001011;
rgb[2898] = 24'b001011000010110100010110;
rgb[2899] = 24'b010000100100010000100010;
rgb[2900] = 24'b010110000101101000101101;
rgb[2901] = 24'b011011100111000100111000;
rgb[2902] = 24'b100001001000100001000100;
rgb[2903] = 24'b100110101001111001001111;
rgb[2904] = 24'b101010111010111101100000;
rgb[2905] = 24'b101101111011101101110110;
rgb[2906] = 24'b110000111100011010001101;
rgb[2907] = 24'b110011111101000110100100;
rgb[2908] = 24'b110110111101110110111011;
rgb[2909] = 24'b111001111110100011010001;
rgb[2910] = 24'b111100111111001111101000;
rgb[2911] = 24'b111111111111111111111111;
rgb[2912] = 24'b000000000000000000000000;
rgb[2913] = 24'b000101110001011100001010;
rgb[2914] = 24'b001011100010111100010100;
rgb[2915] = 24'b010001010100011100011110;
rgb[2916] = 24'b010111000101111100101000;
rgb[2917] = 24'b011100110111011000110011;
rgb[2918] = 24'b100010101000111000111101;
rgb[2919] = 24'b101000101010011001000111;
rgb[2920] = 24'b101100111011011101011000;
rgb[2921] = 24'b101111011100000101110000;
rgb[2922] = 24'b110010001100110010000111;
rgb[2923] = 24'b110100111101011010011111;
rgb[2924] = 24'b110111101110000010110111;
rgb[2925] = 24'b111010011110101011001111;
rgb[2926] = 24'b111101001111010011100111;
rgb[2927] = 24'b111111101111111011111111;
rgb[2928] = 24'b000000000000000000000000;
rgb[2929] = 24'b000110000001100000001001;
rgb[2930] = 24'b001100000011000100010010;
rgb[2931] = 24'b010010000100101000011011;
rgb[2932] = 24'b011000000110001100100100;
rgb[2933] = 24'b011110000111110000101101;
rgb[2934] = 24'b100100011001010100110110;
rgb[2935] = 24'b101010011010111000111111;
rgb[2936] = 24'b101110101011111101010000;
rgb[2937] = 24'b110001001100100001101001;
rgb[2938] = 24'b110011011101000110000010;
rgb[2939] = 24'b110101111101101010011011;
rgb[2940] = 24'b111000011110001110110100;
rgb[2941] = 24'b111010111110110011001101;
rgb[2942] = 24'b111101011111010111100110;
rgb[2943] = 24'b111111111111111111111111;
rgb[2944] = 24'b000000000000000000000000;
rgb[2945] = 24'b000110010001101000000111;
rgb[2946] = 24'b001100100011010000001111;
rgb[2947] = 24'b010010110100111000010111;
rgb[2948] = 24'b011001000110100000011111;
rgb[2949] = 24'b011111101000001000100111;
rgb[2950] = 24'b100101111001110000101111;
rgb[2951] = 24'b101100001011011000110111;
rgb[2952] = 24'b110000011100011101001000;
rgb[2953] = 24'b110010101100111101100010;
rgb[2954] = 24'b110100111101011101111100;
rgb[2955] = 24'b110110111101111110010110;
rgb[2956] = 24'b111001001110011110110000;
rgb[2957] = 24'b111011011110111111001010;
rgb[2958] = 24'b111101101111011111100100;
rgb[2959] = 24'b111111101111111011111111;
rgb[2960] = 24'b000000000000000000000000;
rgb[2961] = 24'b000110100001101100000110;
rgb[2962] = 24'b001101000011011000001101;
rgb[2963] = 24'b010011100101000100010100;
rgb[2964] = 24'b011010000110110000011011;
rgb[2965] = 24'b100000111000100000100001;
rgb[2966] = 24'b100111011010001100101000;
rgb[2967] = 24'b101101111011111000101111;
rgb[2968] = 24'b110010001100111101000000;
rgb[2969] = 24'b110100001101011001011011;
rgb[2970] = 24'b110110001101110101110110;
rgb[2971] = 24'b110111111110001110010010;
rgb[2972] = 24'b111001111110101010101101;
rgb[2973] = 24'b111011111111000111001000;
rgb[2974] = 24'b111101111111100011100011;
rgb[2975] = 24'b111111111111111111111111;
rgb[2976] = 24'b000000000000000000000000;
rgb[2977] = 24'b000110110001110000000101;
rgb[2978] = 24'b001101100011100000001011;
rgb[2979] = 24'b010100010101010100010001;
rgb[2980] = 24'b011011010111000100010110;
rgb[2981] = 24'b100010001000110100011100;
rgb[2982] = 24'b101000111010101000100010;
rgb[2983] = 24'b101111101100011000100111;
rgb[2984] = 24'b110011111101011100111000;
rgb[2985] = 24'b110101101101110101010100;
rgb[2986] = 24'b110111011110001001110001;
rgb[2987] = 24'b111001001110100010001101;
rgb[2988] = 24'b111010101110111010101010;
rgb[2989] = 24'b111100011111001111000110;
rgb[2990] = 24'b111110001111100111100010;
rgb[2991] = 24'b111111101111111011111111;
rgb[2992] = 24'b000000000000000000000000;
rgb[2993] = 24'b000111000001110100000100;
rgb[2994] = 24'b001110000011101000001001;
rgb[2995] = 24'b010101000101100000001101;
rgb[2996] = 24'b011100010111010100010010;
rgb[2997] = 24'b100011011001001100010110;
rgb[2998] = 24'b101010011011000000011011;
rgb[2999] = 24'b110001011100111000011111;
rgb[3000] = 24'b110101101101111100110000;
rgb[3001] = 24'b110111001110001101001110;
rgb[3002] = 24'b111000101110100001101011;
rgb[3003] = 24'b111010001110110010001001;
rgb[3004] = 24'b111011011111000110100110;
rgb[3005] = 24'b111100111111010111000100;
rgb[3006] = 24'b111110011111101011100001;
rgb[3007] = 24'b111111111111111111111111;
rgb[3008] = 24'b000000000000000000000000;
rgb[3009] = 24'b000111010001111000000011;
rgb[3010] = 24'b001110100011110100000110;
rgb[3011] = 24'b010101110101101100001010;
rgb[3012] = 24'b011101010111101000001101;
rgb[3013] = 24'b100100101001100100010000;
rgb[3014] = 24'b101011111011011100010100;
rgb[3015] = 24'b110011011101011000010111;
rgb[3016] = 24'b110111101110011100101000;
rgb[3017] = 24'b111000101110101001000111;
rgb[3018] = 24'b111001111110111001100101;
rgb[3019] = 24'b111011001111000110000100;
rgb[3020] = 24'b111100001111010010100011;
rgb[3021] = 24'b111101011111100011000001;
rgb[3022] = 24'b111110101111101111100000;
rgb[3023] = 24'b111111111111111111111111;
rgb[3024] = 24'b000000000000000000000000;
rgb[3025] = 24'b000111100001111100000010;
rgb[3026] = 24'b001111000011111100000100;
rgb[3027] = 24'b010110100101111100000110;
rgb[3028] = 24'b011110010111111000001001;
rgb[3029] = 24'b100101111001111000001011;
rgb[3030] = 24'b101101011011111000001101;
rgb[3031] = 24'b110101001101111000001111;
rgb[3032] = 24'b111001011110111100100000;
rgb[3033] = 24'b111010001111000101000000;
rgb[3034] = 24'b111011001111001101100000;
rgb[3035] = 24'b111100001111010110000000;
rgb[3036] = 24'b111100111111100010011111;
rgb[3037] = 24'b111101111111101010111111;
rgb[3038] = 24'b111110111111110011011111;
rgb[3039] = 24'b111111111111111111111111;
rgb[3040] = 24'b000000000000000000000000;
rgb[3041] = 24'b000111110010000000000001;
rgb[3042] = 24'b001111100100000100000010;
rgb[3043] = 24'b010111100110001000000011;
rgb[3044] = 24'b011111011000001100000100;
rgb[3045] = 24'b100111001010010000000101;
rgb[3046] = 24'b101111001100010100000110;
rgb[3047] = 24'b110110111110011000000111;
rgb[3048] = 24'b111011001111011100011000;
rgb[3049] = 24'b111011111111100000111001;
rgb[3050] = 24'b111100011111100101011010;
rgb[3051] = 24'b111101001111101001111011;
rgb[3052] = 24'b111101111111101110011100;
rgb[3053] = 24'b111110011111110010111101;
rgb[3054] = 24'b111111001111110111011110;
rgb[3055] = 24'b111111111111111111111111;
rgb[3056] = 24'b000000000000000000000000;
rgb[3057] = 24'b001000000010001000000000;
rgb[3058] = 24'b010000000100010000000000;
rgb[3059] = 24'b011000010110011000000000;
rgb[3060] = 24'b100000011000100000000000;
rgb[3061] = 24'b101000011010101000000000;
rgb[3062] = 24'b110000101100110000000000;
rgb[3063] = 24'b111000101110111000000000;
rgb[3064] = 24'b111100111111111000010001;
rgb[3065] = 24'b111101011111111100110010;
rgb[3066] = 24'b111101101111111001010101;
rgb[3067] = 24'b111110001111111101110110;
rgb[3068] = 24'b111110101111111110011001;
rgb[3069] = 24'b111110111111111110111011;
rgb[3070] = 24'b111111011111111111011101;
rgb[3071] = 24'b111111111111111111111111;
rgb[3072] = 24'b000000000000000000000000;
rgb[3073] = 24'b000100010001000100010001;
rgb[3074] = 24'b001000100010001000100010;
rgb[3075] = 24'b001100110011001100110011;
rgb[3076] = 24'b010001000100010001000100;
rgb[3077] = 24'b010101010101010101010101;
rgb[3078] = 24'b011001100110011001100110;
rgb[3079] = 24'b011101110111011101110111;
rgb[3080] = 24'b100010001000100010001000;
rgb[3081] = 24'b100110011001100110011001;
rgb[3082] = 24'b101010101010101010101010;
rgb[3083] = 24'b101110111011101110111011;
rgb[3084] = 24'b110011001100110011001100;
rgb[3085] = 24'b110111011101110111011101;
rgb[3086] = 24'b111011101110111011101110;
rgb[3087] = 24'b111111111111111111111111;
rgb[3088] = 24'b000000000000000000000000;
rgb[3089] = 24'b000100010001001000001111;
rgb[3090] = 24'b001000110010010000011111;
rgb[3091] = 24'b001101010011011000101111;
rgb[3092] = 24'b010001110100100000111111;
rgb[3093] = 24'b010110010101101001001111;
rgb[3094] = 24'b011010100110110001011111;
rgb[3095] = 24'b011111000111111001101111;
rgb[3096] = 24'b100011011000111110000000;
rgb[3097] = 24'b100111011001111110010010;
rgb[3098] = 24'b101011101010111110100100;
rgb[3099] = 24'b101111101011111110110110;
rgb[3100] = 24'b110011101100111111001000;
rgb[3101] = 24'b110111101101111111011010;
rgb[3102] = 24'b111011101110111111101100;
rgb[3103] = 24'b111111111111111111111111;
rgb[3104] = 24'b000000000000000000000000;
rgb[3105] = 24'b000100100001001100001110;
rgb[3106] = 24'b001001010010011000011101;
rgb[3107] = 24'b001101110011100100101100;
rgb[3108] = 24'b010010100100110100111010;
rgb[3109] = 24'b010111010110000001001001;
rgb[3110] = 24'b011011110111001101011000;
rgb[3111] = 24'b100000101000011001100111;
rgb[3112] = 24'b100100111001011101111000;
rgb[3113] = 24'b101000101010011010001011;
rgb[3114] = 24'b101100101011010110011110;
rgb[3115] = 24'b110000011100010010110001;
rgb[3116] = 24'b110100001101001011000101;
rgb[3117] = 24'b111000001110000111011000;
rgb[3118] = 24'b111011111111000011101011;
rgb[3119] = 24'b111111111111111111111111;
rgb[3120] = 24'b000000000000000000000000;
rgb[3121] = 24'b000100110001010000001101;
rgb[3122] = 24'b001001100010100000011011;
rgb[3123] = 24'b001110100011110100101000;
rgb[3124] = 24'b010011010101000100110110;
rgb[3125] = 24'b011000010110010101000100;
rgb[3126] = 24'b011101000111101001010001;
rgb[3127] = 24'b100010001000111001011111;
rgb[3128] = 24'b100110011001111101110000;
rgb[3129] = 24'b101001111010110110000100;
rgb[3130] = 24'b101101101011101110011000;
rgb[3131] = 24'b110001001100100010101101;
rgb[3132] = 24'b110100111101011011000001;
rgb[3133] = 24'b111000011110001111010110;
rgb[3134] = 24'b111100001111000111101010;
rgb[3135] = 24'b111111111111111111111111;
rgb[3136] = 24'b000000000000000000000000;
rgb[3137] = 24'b000101000001010100001100;
rgb[3138] = 24'b001010000010101100011000;
rgb[3139] = 24'b001111000100000000100101;
rgb[3140] = 24'b010100000101011000110001;
rgb[3141] = 24'b011001010110101100111110;
rgb[3142] = 24'b011110011000000101001010;
rgb[3143] = 24'b100011011001011001010111;
rgb[3144] = 24'b100111101010011101101000;
rgb[3145] = 24'b101011001011010001111101;
rgb[3146] = 24'b101110101100000010010011;
rgb[3147] = 24'b110001111100110110101000;
rgb[3148] = 24'b110101011101100110111110;
rgb[3149] = 24'b111000111110011011010011;
rgb[3150] = 24'b111100011111001011101001;
rgb[3151] = 24'b111111111111111111111111;
rgb[3152] = 24'b000000000000000000000000;
rgb[3153] = 24'b000101010001011000001011;
rgb[3154] = 24'b001010100010110100010110;
rgb[3155] = 24'b001111110100010000100010;
rgb[3156] = 24'b010101000101101000101101;
rgb[3157] = 24'b011010010111000100111000;
rgb[3158] = 24'b011111101000100001000100;
rgb[3159] = 24'b100100111001111001001111;
rgb[3160] = 24'b101001001010111101100000;
rgb[3161] = 24'b101100011011101101110110;
rgb[3162] = 24'b101111101100011010001101;
rgb[3163] = 24'b110010111101000110100100;
rgb[3164] = 24'b110110001101110110111011;
rgb[3165] = 24'b111001011110100011010001;
rgb[3166] = 24'b111100101111001111101000;
rgb[3167] = 24'b111111111111111111111111;
rgb[3168] = 24'b000000000000000000000000;
rgb[3169] = 24'b000101010001011100001010;
rgb[3170] = 24'b001010110010111100010100;
rgb[3171] = 24'b010000010100011100011110;
rgb[3172] = 24'b010101110101111100101000;
rgb[3173] = 24'b011011010111011000110011;
rgb[3174] = 24'b100000111000111000111101;
rgb[3175] = 24'b100110011010011001000111;
rgb[3176] = 24'b101010101011011101011000;
rgb[3177] = 24'b101101101100000101110000;
rgb[3178] = 24'b110000101100110010000111;
rgb[3179] = 24'b110011101101011010011111;
rgb[3180] = 24'b110110101110000010110111;
rgb[3181] = 24'b111001101110101011001111;
rgb[3182] = 24'b111100101111010011100111;
rgb[3183] = 24'b111111101111111011111111;
rgb[3184] = 24'b000000000000000000000000;
rgb[3185] = 24'b000101100001100000001001;
rgb[3186] = 24'b001011010011000100010010;
rgb[3187] = 24'b010001000100101000011011;
rgb[3188] = 24'b010110100110001100100100;
rgb[3189] = 24'b011100010111110000101101;
rgb[3190] = 24'b100010001001010100110110;
rgb[3191] = 24'b100111101010111000111111;
rgb[3192] = 24'b101011111011111101010000;
rgb[3193] = 24'b101110111100100001101001;
rgb[3194] = 24'b110001101101000110000010;
rgb[3195] = 24'b110100011101101010011011;
rgb[3196] = 24'b110111011110001110110100;
rgb[3197] = 24'b111010001110110011001101;
rgb[3198] = 24'b111100111111010111100110;
rgb[3199] = 24'b111111111111111111111111;
rgb[3200] = 24'b000000000000000000000000;
rgb[3201] = 24'b000101110001101000000111;
rgb[3202] = 24'b001011100011010000001111;
rgb[3203] = 24'b010001100100111000010111;
rgb[3204] = 24'b010111010110100000011111;
rgb[3205] = 24'b011101011000001000100111;
rgb[3206] = 24'b100011001001110000101111;
rgb[3207] = 24'b101001001011011000110111;
rgb[3208] = 24'b101101011100011101001000;
rgb[3209] = 24'b101111111100111101100010;
rgb[3210] = 24'b110010101101011101111100;
rgb[3211] = 24'b110101001101111110010110;
rgb[3212] = 24'b110111111110011110110000;
rgb[3213] = 24'b111010011110111111001010;
rgb[3214] = 24'b111101001111011111100100;
rgb[3215] = 24'b111111101111111011111111;
rgb[3216] = 24'b000000000000000000000000;
rgb[3217] = 24'b000110000001101100000110;
rgb[3218] = 24'b001100000011011000001101;
rgb[3219] = 24'b010010000101000100010100;
rgb[3220] = 24'b011000010110110000011011;
rgb[3221] = 24'b011110011000100000100001;
rgb[3222] = 24'b100100011010001100101000;
rgb[3223] = 24'b101010101011111000101111;
rgb[3224] = 24'b101110111100111101000000;
rgb[3225] = 24'b110001001101011001011011;
rgb[3226] = 24'b110011101101110101110110;
rgb[3227] = 24'b110110001110001110010010;
rgb[3228] = 24'b111000011110101010101101;
rgb[3229] = 24'b111010111111000111001000;
rgb[3230] = 24'b111101011111100011100011;
rgb[3231] = 24'b111111111111111111111111;
rgb[3232] = 24'b000000000000000000000000;
rgb[3233] = 24'b000110010001110000000101;
rgb[3234] = 24'b001100100011100000001011;
rgb[3235] = 24'b010010110101010100010001;
rgb[3236] = 24'b011001000111000100010110;
rgb[3237] = 24'b011111011000110100011100;
rgb[3238] = 24'b100101101010101000100010;
rgb[3239] = 24'b101011111100011000100111;
rgb[3240] = 24'b110000001101011100111000;
rgb[3241] = 24'b110010011101110101010100;
rgb[3242] = 24'b110100101110001001110001;
rgb[3243] = 24'b110110111110100010001101;
rgb[3244] = 24'b111001001110111010101010;
rgb[3245] = 24'b111011011111001111000110;
rgb[3246] = 24'b111101101111100111100010;
rgb[3247] = 24'b111111101111111011111111;
rgb[3248] = 24'b000000000000000000000000;
rgb[3249] = 24'b000110010001110100000100;
rgb[3250] = 24'b001100110011101000001001;
rgb[3251] = 24'b010011010101100000001101;
rgb[3252] = 24'b011001110111010100010010;
rgb[3253] = 24'b100000011001001100010110;
rgb[3254] = 24'b100110111011000000011011;
rgb[3255] = 24'b101101011100111000011111;
rgb[3256] = 24'b110001101101111100110000;
rgb[3257] = 24'b110011101110001101001110;
rgb[3258] = 24'b110101101110100001101011;
rgb[3259] = 24'b110111101110110010001001;
rgb[3260] = 24'b111001101111000110100110;
rgb[3261] = 24'b111011101111010111000100;
rgb[3262] = 24'b111101101111101011100001;
rgb[3263] = 24'b111111111111111111111111;
rgb[3264] = 24'b000000000000000000000000;
rgb[3265] = 24'b000110100001111000000011;
rgb[3266] = 24'b001101010011110100000110;
rgb[3267] = 24'b010100000101101100001010;
rgb[3268] = 24'b011010100111101000001101;
rgb[3269] = 24'b100001011001100100010000;
rgb[3270] = 24'b101000001011011100010100;
rgb[3271] = 24'b101110111101011000010111;
rgb[3272] = 24'b110011001110011100101000;
rgb[3273] = 24'b110100111110101001000111;
rgb[3274] = 24'b110110101110111001100101;
rgb[3275] = 24'b111000011111000110000100;
rgb[3276] = 24'b111010011111010010100011;
rgb[3277] = 24'b111100001111100011000001;
rgb[3278] = 24'b111101111111101111100000;
rgb[3279] = 24'b111111111111111111111111;
rgb[3280] = 24'b000000000000000000000000;
rgb[3281] = 24'b000110110001111100000010;
rgb[3282] = 24'b001101110011111100000100;
rgb[3283] = 24'b010100100101111100000110;
rgb[3284] = 24'b011011100111111000001001;
rgb[3285] = 24'b100010011001111000001011;
rgb[3286] = 24'b101001011011111000001101;
rgb[3287] = 24'b110000001101111000001111;
rgb[3288] = 24'b110100011110111100100000;
rgb[3289] = 24'b110110001111000101000000;
rgb[3290] = 24'b110111101111001101100000;
rgb[3291] = 24'b111001011111010110000000;
rgb[3292] = 24'b111010111111100010011111;
rgb[3293] = 24'b111100101111101010111111;
rgb[3294] = 24'b111110001111110011011111;
rgb[3295] = 24'b111111111111111111111111;
rgb[3296] = 24'b000000000000000000000000;
rgb[3297] = 24'b000111000010000000000001;
rgb[3298] = 24'b001110000100000100000010;
rgb[3299] = 24'b010101010110001000000011;
rgb[3300] = 24'b011100011000001100000100;
rgb[3301] = 24'b100011011010010000000101;
rgb[3302] = 24'b101010101100010100000110;
rgb[3303] = 24'b110001101110011000000111;
rgb[3304] = 24'b110101111111011100011000;
rgb[3305] = 24'b110111011111100000111001;
rgb[3306] = 24'b111000101111100101011010;
rgb[3307] = 24'b111010001111101001111011;
rgb[3308] = 24'b111011101111101110011100;
rgb[3309] = 24'b111100111111110010111101;
rgb[3310] = 24'b111110011111110111011110;
rgb[3311] = 24'b111111111111111111111111;
rgb[3312] = 24'b000000000000000000000000;
rgb[3313] = 24'b000111010010001000000000;
rgb[3314] = 24'b001110100100010000000000;
rgb[3315] = 24'b010101110110011000000000;
rgb[3316] = 24'b011101001000100000000000;
rgb[3317] = 24'b100100011010101000000000;
rgb[3318] = 24'b101011101100110000000000;
rgb[3319] = 24'b110011001110111000000000;
rgb[3320] = 24'b110111011111111000010001;
rgb[3321] = 24'b111000011111111100110010;
rgb[3322] = 24'b111001101111111001010101;
rgb[3323] = 24'b111010111111111101110110;
rgb[3324] = 24'b111100001111111110011001;
rgb[3325] = 24'b111101011111111110111011;
rgb[3326] = 24'b111110101111111111011101;
rgb[3327] = 24'b111111111111111111111111;
rgb[3328] = 24'b000000000000000000000000;
rgb[3329] = 24'b000100010001000100010001;
rgb[3330] = 24'b001000100010001000100010;
rgb[3331] = 24'b001100110011001100110011;
rgb[3332] = 24'b010001000100010001000100;
rgb[3333] = 24'b010101010101010101010101;
rgb[3334] = 24'b011001100110011001100110;
rgb[3335] = 24'b011101110111011101110111;
rgb[3336] = 24'b100010001000100010001000;
rgb[3337] = 24'b100110011001100110011001;
rgb[3338] = 24'b101010101010101010101010;
rgb[3339] = 24'b101110111011101110111011;
rgb[3340] = 24'b110011001100110011001100;
rgb[3341] = 24'b110111011101110111011101;
rgb[3342] = 24'b111011101110111011101110;
rgb[3343] = 24'b111111111111111111111111;
rgb[3344] = 24'b000000000000000000000000;
rgb[3345] = 24'b000100010001001000001111;
rgb[3346] = 24'b001000110010010000011111;
rgb[3347] = 24'b001101000011011000101111;
rgb[3348] = 24'b010001100100100000111111;
rgb[3349] = 24'b010101110101101001001111;
rgb[3350] = 24'b011010010110110001011111;
rgb[3351] = 24'b011110110111111001101111;
rgb[3352] = 24'b100011001000111110000000;
rgb[3353] = 24'b100111001001111110010010;
rgb[3354] = 24'b101011001010111110100100;
rgb[3355] = 24'b101111011011111110110110;
rgb[3356] = 24'b110011011100111111001000;
rgb[3357] = 24'b110111101101111111011010;
rgb[3358] = 24'b111011101110111111101100;
rgb[3359] = 24'b111111111111111111111111;
rgb[3360] = 24'b000000000000000000000000;
rgb[3361] = 24'b000100100001001100001110;
rgb[3362] = 24'b001001000010011000011101;
rgb[3363] = 24'b001101100011100100101100;
rgb[3364] = 24'b010010000100110100111010;
rgb[3365] = 24'b010110100110000001001001;
rgb[3366] = 24'b011011010111001101011000;
rgb[3367] = 24'b011111111000011001100111;
rgb[3368] = 24'b100100001001011101111000;
rgb[3369] = 24'b101000001010011010001011;
rgb[3370] = 24'b101011111011010110011110;
rgb[3371] = 24'b101111111100010010110001;
rgb[3372] = 24'b110011111101001011000101;
rgb[3373] = 24'b110111111110000111011000;
rgb[3374] = 24'b111011111111000011101011;
rgb[3375] = 24'b111111111111111111111111;
rgb[3376] = 24'b000000000000000000000000;
rgb[3377] = 24'b000100100001010000001101;
rgb[3378] = 24'b001001010010100000011011;
rgb[3379] = 24'b001110000011110100101000;
rgb[3380] = 24'b010010110101000100110110;
rgb[3381] = 24'b010111010110010101000100;
rgb[3382] = 24'b011100000111101001010001;
rgb[3383] = 24'b100000111000111001011111;
rgb[3384] = 24'b100101001001111101110000;
rgb[3385] = 24'b101000111010110110000100;
rgb[3386] = 24'b101100101011101110011000;
rgb[3387] = 24'b110000101100100010101101;
rgb[3388] = 24'b110100011101011011000001;
rgb[3389] = 24'b111000001110001111010110;
rgb[3390] = 24'b111011111111000111101010;
rgb[3391] = 24'b111111111111111111111111;
rgb[3392] = 24'b000000000000000000000000;
rgb[3393] = 24'b000100110001010100001100;
rgb[3394] = 24'b001001100010101100011000;
rgb[3395] = 24'b001110100100000000100101;
rgb[3396] = 24'b010011010101011000110001;
rgb[3397] = 24'b011000000110101100111110;
rgb[3398] = 24'b011101001000000101001010;
rgb[3399] = 24'b100001111001011001010111;
rgb[3400] = 24'b100110001010011101101000;
rgb[3401] = 24'b101001111011010001111101;
rgb[3402] = 24'b101101011100000010010011;
rgb[3403] = 24'b110001001100110110101000;
rgb[3404] = 24'b110100111101100110111110;
rgb[3405] = 24'b111000011110011011010011;
rgb[3406] = 24'b111100001111001011101001;
rgb[3407] = 24'b111111111111111111111111;
rgb[3408] = 24'b000000000000000000000000;
rgb[3409] = 24'b000100110001011000001011;
rgb[3410] = 24'b001001110010110100010110;
rgb[3411] = 24'b001110110100010000100010;
rgb[3412] = 24'b010011110101101000101101;
rgb[3413] = 24'b011000110111000100111000;
rgb[3414] = 24'b011101111000100001000100;
rgb[3415] = 24'b100010111001111001001111;
rgb[3416] = 24'b100111001010111101100000;
rgb[3417] = 24'b101010101011101101110110;
rgb[3418] = 24'b101110001100011010001101;
rgb[3419] = 24'b110001101101000110100100;
rgb[3420] = 24'b110101001101110110111011;
rgb[3421] = 24'b111000101110100011010001;
rgb[3422] = 24'b111100001111001111101000;
rgb[3423] = 24'b111111111111111111111111;
rgb[3424] = 24'b000000000000000000000000;
rgb[3425] = 24'b000101000001011100001010;
rgb[3426] = 24'b001010010010111100010100;
rgb[3427] = 24'b001111010100011100011110;
rgb[3428] = 24'b010100100101111100101000;
rgb[3429] = 24'b011001100111011000110011;
rgb[3430] = 24'b011110111000111000111101;
rgb[3431] = 24'b100011111010011001000111;
rgb[3432] = 24'b101000001011011101011000;
rgb[3433] = 24'b101011101100000101110000;
rgb[3434] = 24'b101110111100110010000111;
rgb[3435] = 24'b110010011101011010011111;
rgb[3436] = 24'b110101101110000010110111;
rgb[3437] = 24'b111001001110101011001111;
rgb[3438] = 24'b111100011111010011100111;
rgb[3439] = 24'b111111101111111011111111;
rgb[3440] = 24'b000000000000000000000000;
rgb[3441] = 24'b000101010001100000001001;
rgb[3442] = 24'b001010100011000100010010;
rgb[3443] = 24'b001111110100101000011011;
rgb[3444] = 24'b010101000110001100100100;
rgb[3445] = 24'b011010010111110000101101;
rgb[3446] = 24'b011111101001010100110110;
rgb[3447] = 24'b100101001010111000111111;
rgb[3448] = 24'b101001011011111101010000;
rgb[3449] = 24'b101100011100100001101001;
rgb[3450] = 24'b101111101101000110000010;
rgb[3451] = 24'b110010111101101010011011;
rgb[3452] = 24'b110110001110001110110100;
rgb[3453] = 24'b111001011110110011001101;
rgb[3454] = 24'b111100101111010111100110;
rgb[3455] = 24'b111111111111111111111111;
rgb[3456] = 24'b000000000000000000000000;
rgb[3457] = 24'b000101010001101000000111;
rgb[3458] = 24'b001010110011010000001111;
rgb[3459] = 24'b010000010100111000010111;
rgb[3460] = 24'b010101100110100000011111;
rgb[3461] = 24'b011011001000001000100111;
rgb[3462] = 24'b100000101001110000101111;
rgb[3463] = 24'b100110001011011000110111;
rgb[3464] = 24'b101010011100011101001000;
rgb[3465] = 24'b101101011100111101100010;
rgb[3466] = 24'b110000011101011101111100;
rgb[3467] = 24'b110011011101111110010110;
rgb[3468] = 24'b110110101110011110110000;
rgb[3469] = 24'b111001101110111111001010;
rgb[3470] = 24'b111100101111011111100100;
rgb[3471] = 24'b111111101111111011111111;
rgb[3472] = 24'b000000000000000000000000;
rgb[3473] = 24'b000101100001101100000110;
rgb[3474] = 24'b001011000011011000001101;
rgb[3475] = 24'b010000110101000100010100;
rgb[3476] = 24'b010110010110110000011011;
rgb[3477] = 24'b011011111000100000100001;
rgb[3478] = 24'b100001101010001100101000;
rgb[3479] = 24'b100111001011111000101111;
rgb[3480] = 24'b101011011100111101000000;
rgb[3481] = 24'b101110011101011001011011;
rgb[3482] = 24'b110001001101110101110110;
rgb[3483] = 24'b110100001110001110010010;
rgb[3484] = 24'b110111001110101010101101;
rgb[3485] = 24'b111001111111000111001000;
rgb[3486] = 24'b111100111111100011100011;
rgb[3487] = 24'b111111111111111111111111;
rgb[3488] = 24'b000000000000000000000000;
rgb[3489] = 24'b000101100001110000000101;
rgb[3490] = 24'b001011010011100000001011;
rgb[3491] = 24'b010001000101010100010001;
rgb[3492] = 24'b010110110111000100010110;
rgb[3493] = 24'b011100101000110100011100;
rgb[3494] = 24'b100010011010101000100010;
rgb[3495] = 24'b101000001100011000100111;
rgb[3496] = 24'b101100011101011100111000;
rgb[3497] = 24'b101111001101110101010100;
rgb[3498] = 24'b110001111110001001110001;
rgb[3499] = 24'b110100101110100010001101;
rgb[3500] = 24'b110111011110111010101010;
rgb[3501] = 24'b111010001111001111000110;
rgb[3502] = 24'b111100111111100111100010;
rgb[3503] = 24'b111111101111111011111111;
rgb[3504] = 24'b000000000000000000000000;
rgb[3505] = 24'b000101110001110100000100;
rgb[3506] = 24'b001011110011101000001001;
rgb[3507] = 24'b010001100101100000001101;
rgb[3508] = 24'b010111100111010100010010;
rgb[3509] = 24'b011101011001001100010110;
rgb[3510] = 24'b100011011011000000011011;
rgb[3511] = 24'b101001001100111000011111;
rgb[3512] = 24'b101101011101111100110000;
rgb[3513] = 24'b110000001110001101001110;
rgb[3514] = 24'b110010101110100001101011;
rgb[3515] = 24'b110101011110110010001001;
rgb[3516] = 24'b110111111111000110100110;
rgb[3517] = 24'b111010101111010111000100;
rgb[3518] = 24'b111101001111101011100001;
rgb[3519] = 24'b111111111111111111111111;
rgb[3520] = 24'b000000000000000000000000;
rgb[3521] = 24'b000110000001111000000011;
rgb[3522] = 24'b001100000011110100000110;
rgb[3523] = 24'b010010000101101100001010;
rgb[3524] = 24'b011000000111101000001101;
rgb[3525] = 24'b011110001001100100010000;
rgb[3526] = 24'b100100001011011100010100;
rgb[3527] = 24'b101010001101011000010111;
rgb[3528] = 24'b101110011110011100101000;
rgb[3529] = 24'b110000111110101001000111;
rgb[3530] = 24'b110011011110111001100101;
rgb[3531] = 24'b110101111111000110000100;
rgb[3532] = 24'b111000011111010010100011;
rgb[3533] = 24'b111010111111100011000001;
rgb[3534] = 24'b111101011111101111100000;
rgb[3535] = 24'b111111111111111111111111;
rgb[3536] = 24'b000000000000000000000000;
rgb[3537] = 24'b000110000001111100000010;
rgb[3538] = 24'b001100010011111100000100;
rgb[3539] = 24'b010010100101111100000110;
rgb[3540] = 24'b011000100111111000001001;
rgb[3541] = 24'b011110111001111000001011;
rgb[3542] = 24'b100101001011111000001101;
rgb[3543] = 24'b101011011101111000001111;
rgb[3544] = 24'b101111101110111100100000;
rgb[3545] = 24'b110001111111000101000000;
rgb[3546] = 24'b110100001111001101100000;
rgb[3547] = 24'b110110011111010110000000;
rgb[3548] = 24'b111000111111100010011111;
rgb[3549] = 24'b111011001111101010111111;
rgb[3550] = 24'b111101011111110011011111;
rgb[3551] = 24'b111111111111111111111111;
rgb[3552] = 24'b000000000000000000000000;
rgb[3553] = 24'b000110010010000000000001;
rgb[3554] = 24'b001100100100000100000010;
rgb[3555] = 24'b010010110110001000000011;
rgb[3556] = 24'b011001011000001100000100;
rgb[3557] = 24'b011111101010010000000101;
rgb[3558] = 24'b100101111100010100000110;
rgb[3559] = 24'b101100011110011000000111;
rgb[3560] = 24'b110000101111011100011000;
rgb[3561] = 24'b110010101111100000111001;
rgb[3562] = 24'b110100111111100101011010;
rgb[3563] = 24'b110111001111101001111011;
rgb[3564] = 24'b111001001111101110011100;
rgb[3565] = 24'b111011011111110010111101;
rgb[3566] = 24'b111101101111110111011110;
rgb[3567] = 24'b111111111111111111111111;
rgb[3568] = 24'b000000000000000000000000;
rgb[3569] = 24'b000110010010001000000000;
rgb[3570] = 24'b001100110100010000000000;
rgb[3571] = 24'b010011010110011000000000;
rgb[3572] = 24'b011001111000100000000000;
rgb[3573] = 24'b100000011010101000000000;
rgb[3574] = 24'b100110111100110000000000;
rgb[3575] = 24'b101101011110111000000000;
rgb[3576] = 24'b110001101111111000010001;
rgb[3577] = 24'b110011101111111100110010;
rgb[3578] = 24'b110101101111111001010101;
rgb[3579] = 24'b110111101111111101110110;
rgb[3580] = 24'b111001101111111110011001;
rgb[3581] = 24'b111011101111111110111011;
rgb[3582] = 24'b111101101111111111011101;
rgb[3583] = 24'b111111111111111111111111;
rgb[3584] = 24'b000000000000000000000000;
rgb[3585] = 24'b000100010001000100010001;
rgb[3586] = 24'b001000100010001000100010;
rgb[3587] = 24'b001100110011001100110011;
rgb[3588] = 24'b010001000100010001000100;
rgb[3589] = 24'b010101010101010101010101;
rgb[3590] = 24'b011001100110011001100110;
rgb[3591] = 24'b011101110111011101110111;
rgb[3592] = 24'b100010001000100010001000;
rgb[3593] = 24'b100110011001100110011001;
rgb[3594] = 24'b101010101010101010101010;
rgb[3595] = 24'b101110111011101110111011;
rgb[3596] = 24'b110011001100110011001100;
rgb[3597] = 24'b110111011101110111011101;
rgb[3598] = 24'b111011101110111011101110;
rgb[3599] = 24'b111111111111111111111111;
rgb[3600] = 24'b000000000000000000000000;
rgb[3601] = 24'b000100010001001000001111;
rgb[3602] = 24'b001000100010010000011111;
rgb[3603] = 24'b001101000011011000101111;
rgb[3604] = 24'b010001010100100000111111;
rgb[3605] = 24'b010101100101101001001111;
rgb[3606] = 24'b011010000110110001011111;
rgb[3607] = 24'b011110010111111001101111;
rgb[3608] = 24'b100010101000111110000000;
rgb[3609] = 24'b100110111001111110010010;
rgb[3610] = 24'b101010111010111110100100;
rgb[3611] = 24'b101111001011111110110110;
rgb[3612] = 24'b110011011100111111001000;
rgb[3613] = 24'b110111011101111111011010;
rgb[3614] = 24'b111011101110111111101100;
rgb[3615] = 24'b111111111111111111111111;
rgb[3616] = 24'b000000000000000000000000;
rgb[3617] = 24'b000100010001001100001110;
rgb[3618] = 24'b001000110010011000011101;
rgb[3619] = 24'b001101010011100100101100;
rgb[3620] = 24'b010001110100110100111010;
rgb[3621] = 24'b010110000110000001001001;
rgb[3622] = 24'b011010100111001101011000;
rgb[3623] = 24'b011111001000011001100111;
rgb[3624] = 24'b100011011001011101111000;
rgb[3625] = 24'b100111011010011010001011;
rgb[3626] = 24'b101011011011010110011110;
rgb[3627] = 24'b101111101100010010110001;
rgb[3628] = 24'b110011101101001011000101;
rgb[3629] = 24'b110111101110000111011000;
rgb[3630] = 24'b111011101111000011101011;
rgb[3631] = 24'b111111111111111111111111;
rgb[3632] = 24'b000000000000000000000000;
rgb[3633] = 24'b000100100001010000001101;
rgb[3634] = 24'b001001000010100000011011;
rgb[3635] = 24'b001101100011110100101000;
rgb[3636] = 24'b010010000101000100110110;
rgb[3637] = 24'b010110100110010101000100;
rgb[3638] = 24'b011011000111101001010001;
rgb[3639] = 24'b011111101000111001011111;
rgb[3640] = 24'b100011111001111101110000;
rgb[3641] = 24'b100111111010110110000100;
rgb[3642] = 24'b101011111011101110011000;
rgb[3643] = 24'b101111111100100010101101;
rgb[3644] = 24'b110011111101011011000001;
rgb[3645] = 24'b110111111110001111010110;
rgb[3646] = 24'b111011111111000111101010;
rgb[3647] = 24'b111111111111111111111111;
rgb[3648] = 24'b000000000000000000000000;
rgb[3649] = 24'b000100100001010100001100;
rgb[3650] = 24'b001001010010101100011000;
rgb[3651] = 24'b001101110100000000100101;
rgb[3652] = 24'b010010100101011000110001;
rgb[3653] = 24'b010111000110101100111110;
rgb[3654] = 24'b011011111000000101001010;
rgb[3655] = 24'b100000011001011001010111;
rgb[3656] = 24'b100100101010011101101000;
rgb[3657] = 24'b101000101011010001111101;
rgb[3658] = 24'b101100011100000010010011;
rgb[3659] = 24'b110000011100110110101000;
rgb[3660] = 24'b110100001101100110111110;
rgb[3661] = 24'b111000001110011011010011;
rgb[3662] = 24'b111011111111001011101001;
rgb[3663] = 24'b111111111111111111111111;
rgb[3664] = 24'b000000000000000000000000;
rgb[3665] = 24'b000100100001011000001011;
rgb[3666] = 24'b001001010010110100010110;
rgb[3667] = 24'b001110000100010000100010;
rgb[3668] = 24'b010010110101101000101101;
rgb[3669] = 24'b010111100111000100111000;
rgb[3670] = 24'b011100011000100001000100;
rgb[3671] = 24'b100001001001111001001111;
rgb[3672] = 24'b100101011010111101100000;
rgb[3673] = 24'b101001001011101101110110;
rgb[3674] = 24'b101100111100011010001101;
rgb[3675] = 24'b110000101101000110100100;
rgb[3676] = 24'b110100011101110110111011;
rgb[3677] = 24'b111000001110100011010001;
rgb[3678] = 24'b111011111111001111101000;
rgb[3679] = 24'b111111111111111111111111;
rgb[3680] = 24'b000000000000000000000000;
rgb[3681] = 24'b000100110001011100001010;
rgb[3682] = 24'b001001100010111100010100;
rgb[3683] = 24'b001110010100011100011110;
rgb[3684] = 24'b010011010101111100101000;
rgb[3685] = 24'b011000000111011000110011;
rgb[3686] = 24'b011100111000111000111101;
rgb[3687] = 24'b100001101010011001000111;
rgb[3688] = 24'b100101111011011101011000;
rgb[3689] = 24'b101001101100000101110000;
rgb[3690] = 24'b101101011100110010000111;
rgb[3691] = 24'b110001001101011010011111;
rgb[3692] = 24'b110100101110000010110111;
rgb[3693] = 24'b111000011110101011001111;
rgb[3694] = 24'b111100001111010011100111;
rgb[3695] = 24'b111111101111111011111111;
rgb[3696] = 24'b000000000000000000000000;
rgb[3697] = 24'b000100110001100000001001;
rgb[3698] = 24'b001001110011000100010010;
rgb[3699] = 24'b001110100100101000011011;
rgb[3700] = 24'b010011100110001100100100;
rgb[3701] = 24'b011000100111110000101101;
rgb[3702] = 24'b011101011001010100110110;
rgb[3703] = 24'b100010011010111000111111;
rgb[3704] = 24'b100110101011111101010000;
rgb[3705] = 24'b101010001100100001101001;
rgb[3706] = 24'b101101111101000110000010;
rgb[3707] = 24'b110001011101101010011011;
rgb[3708] = 24'b110100111110001110110100;
rgb[3709] = 24'b111000101110110011001101;
rgb[3710] = 24'b111100001111010111100110;
rgb[3711] = 24'b111111111111111111111111;
rgb[3712] = 24'b000000000000000000000000;
rgb[3713] = 24'b000101000001101000000111;
rgb[3714] = 24'b001010000011010000001111;
rgb[3715] = 24'b001111000100111000010111;
rgb[3716] = 24'b010100000110100000011111;
rgb[3717] = 24'b011001001000001000100111;
rgb[3718] = 24'b011110001001110000101111;
rgb[3719] = 24'b100011001011011000110111;
rgb[3720] = 24'b100111011100011101001000;
rgb[3721] = 24'b101010111100111101100010;
rgb[3722] = 24'b101110011101011101111100;
rgb[3723] = 24'b110001111101111110010110;
rgb[3724] = 24'b110101011110011110110000;
rgb[3725] = 24'b111000111110111111001010;
rgb[3726] = 24'b111100011111011111100100;
rgb[3727] = 24'b111111101111111011111111;
rgb[3728] = 24'b000000000000000000000000;
rgb[3729] = 24'b000101000001101100000110;
rgb[3730] = 24'b001010000011011000001101;
rgb[3731] = 24'b001111010101000100010100;
rgb[3732] = 24'b010100010110110000011011;
rgb[3733] = 24'b011001011000100000100001;
rgb[3734] = 24'b011110101010001100101000;
rgb[3735] = 24'b100011101011111000101111;
rgb[3736] = 24'b100111111100111101000000;
rgb[3737] = 24'b101011011101011001011011;
rgb[3738] = 24'b101110101101110101110110;
rgb[3739] = 24'b110010001110001110010010;
rgb[3740] = 24'b110101101110101010101101;
rgb[3741] = 24'b111000111111000111001000;
rgb[3742] = 24'b111100011111100011100011;
rgb[3743] = 24'b111111111111111111111111;
rgb[3744] = 24'b000000000000000000000000;
rgb[3745] = 24'b000101000001110000000101;
rgb[3746] = 24'b001010010011100000001011;
rgb[3747] = 24'b001111100101010100010001;
rgb[3748] = 24'b010100110111000100010110;
rgb[3749] = 24'b011001111000110100011100;
rgb[3750] = 24'b011111001010101000100010;
rgb[3751] = 24'b100100011100011000100111;
rgb[3752] = 24'b101000101101011100111000;
rgb[3753] = 24'b101011111101110101010100;
rgb[3754] = 24'b101111001110001001110001;
rgb[3755] = 24'b110010101110100010001101;
rgb[3756] = 24'b110101111110111010101010;
rgb[3757] = 24'b111001001111001111000110;
rgb[3758] = 24'b111100011111100111100010;
rgb[3759] = 24'b111111101111111011111111;
rgb[3760] = 24'b000000000000000000000000;
rgb[3761] = 24'b000101010001110100000100;
rgb[3762] = 24'b001010100011101000001001;
rgb[3763] = 24'b001111110101100000001101;
rgb[3764] = 24'b010101000111010100010010;
rgb[3765] = 24'b011010011001001100010110;
rgb[3766] = 24'b011111101011000000011011;
rgb[3767] = 24'b100101001100111000011111;
rgb[3768] = 24'b101001011101111100110000;
rgb[3769] = 24'b101100011110001101001110;
rgb[3770] = 24'b101111101110100001101011;
rgb[3771] = 24'b110010111110110010001001;
rgb[3772] = 24'b110110001111000110100110;
rgb[3773] = 24'b111001011111010111000100;
rgb[3774] = 24'b111100101111101011100001;
rgb[3775] = 24'b111111111111111111111111;
rgb[3776] = 24'b000000000000000000000000;
rgb[3777] = 24'b000101010001111000000011;
rgb[3778] = 24'b001010110011110100000110;
rgb[3779] = 24'b010000000101101100001010;
rgb[3780] = 24'b010101100111101000001101;
rgb[3781] = 24'b011010111001100100010000;
rgb[3782] = 24'b100000011011011100010100;
rgb[3783] = 24'b100101101101011000010111;
rgb[3784] = 24'b101001111110011100101000;
rgb[3785] = 24'b101101001110101001000111;
rgb[3786] = 24'b110000001110111001100101;
rgb[3787] = 24'b110011011111000110000100;
rgb[3788] = 24'b110110011111010010100011;
rgb[3789] = 24'b111001101111100011000001;
rgb[3790] = 24'b111100101111101111100000;
rgb[3791] = 24'b111111111111111111111111;
rgb[3792] = 24'b000000000000000000000000;
rgb[3793] = 24'b000101010001111100000010;
rgb[3794] = 24'b001010110011111100000100;
rgb[3795] = 24'b010000010101111100000110;
rgb[3796] = 24'b010101110111111000001001;
rgb[3797] = 24'b011011011001111000001011;
rgb[3798] = 24'b100000111011111000001101;
rgb[3799] = 24'b100110011101111000001111;
rgb[3800] = 24'b101010101110111100100000;
rgb[3801] = 24'b101101101111000101000000;
rgb[3802] = 24'b110000101111001101100000;
rgb[3803] = 24'b110011101111010110000000;
rgb[3804] = 24'b110110101111100010011111;
rgb[3805] = 24'b111001101111101010111111;
rgb[3806] = 24'b111100101111110011011111;
rgb[3807] = 24'b111111111111111111111111;
rgb[3808] = 24'b000000000000000000000000;
rgb[3809] = 24'b000101100010000000000001;
rgb[3810] = 24'b001011000100000100000010;
rgb[3811] = 24'b010000100110001000000011;
rgb[3812] = 24'b010110011000001100000100;
rgb[3813] = 24'b011011111010010000000101;
rgb[3814] = 24'b100001011100010100000110;
rgb[3815] = 24'b100111001110011000000111;
rgb[3816] = 24'b101011011111011100011000;
rgb[3817] = 24'b101110001111100000111001;
rgb[3818] = 24'b110001001111100101011010;
rgb[3819] = 24'b110100001111101001111011;
rgb[3820] = 24'b110110111111101110011100;
rgb[3821] = 24'b111001111111110010111101;
rgb[3822] = 24'b111100111111110111011110;
rgb[3823] = 24'b111111111111111111111111;
rgb[3824] = 24'b000000000000000000000000;
rgb[3825] = 24'b000101100010001000000000;
rgb[3826] = 24'b001011010100010000000000;
rgb[3827] = 24'b010000110110011000000000;
rgb[3828] = 24'b010110101000100000000000;
rgb[3829] = 24'b011100011010101000000000;
rgb[3830] = 24'b100001111100110000000000;
rgb[3831] = 24'b100111101110111000000000;
rgb[3832] = 24'b101011111111111000010001;
rgb[3833] = 24'b101110101111111100110010;
rgb[3834] = 24'b110001101111111001010101;
rgb[3835] = 24'b110100011111111101110110;
rgb[3836] = 24'b110111001111111110011001;
rgb[3837] = 24'b111010001111111110111011;
rgb[3838] = 24'b111100111111111111011101;
rgb[3839] = 24'b111111111111111111111111;
rgb[3840] = 24'b000000000000000000000000;
rgb[3841] = 24'b000100010001000100010001;
rgb[3842] = 24'b001000100010001000100010;
rgb[3843] = 24'b001100110011001100110011;
rgb[3844] = 24'b010001000100010001000100;
rgb[3845] = 24'b010101010101010101010101;
rgb[3846] = 24'b011001100110011001100110;
rgb[3847] = 24'b011101110111011101110111;
rgb[3848] = 24'b100010001000100010001000;
rgb[3849] = 24'b100110011001100110011001;
rgb[3850] = 24'b101010101010101010101010;
rgb[3851] = 24'b101110111011101110111011;
rgb[3852] = 24'b110011001100110011001100;
rgb[3853] = 24'b110111011101110111011101;
rgb[3854] = 24'b111011101110111011101110;
rgb[3855] = 24'b111111111111111111111111;
rgb[3856] = 24'b000000000000000000000000;
rgb[3857] = 24'b000100010001001000001111;
rgb[3858] = 24'b001000100010010000011111;
rgb[3859] = 24'b001100110011011000101111;
rgb[3860] = 24'b010001000100100000111111;
rgb[3861] = 24'b010101010101101001001111;
rgb[3862] = 24'b011001100110110001011111;
rgb[3863] = 24'b011110000111111001101111;
rgb[3864] = 24'b100010011000111110000000;
rgb[3865] = 24'b100110011001111110010010;
rgb[3866] = 24'b101010101010111110100100;
rgb[3867] = 24'b101110111011111110110110;
rgb[3868] = 24'b110011001100111111001000;
rgb[3869] = 24'b110111011101111111011010;
rgb[3870] = 24'b111011101110111111101100;
rgb[3871] = 24'b111111111111111111111111;
rgb[3872] = 24'b000000000000000000000000;
rgb[3873] = 24'b000100010001001100001110;
rgb[3874] = 24'b001000100010011000011101;
rgb[3875] = 24'b001100110011100100101100;
rgb[3876] = 24'b010001010100110100111010;
rgb[3877] = 24'b010101100110000001001001;
rgb[3878] = 24'b011001110111001101011000;
rgb[3879] = 24'b011110011000011001100111;
rgb[3880] = 24'b100010101001011101111000;
rgb[3881] = 24'b100110101010011010001011;
rgb[3882] = 24'b101010111011010110011110;
rgb[3883] = 24'b101111001100010010110001;
rgb[3884] = 24'b110011001101001011000101;
rgb[3885] = 24'b110111011110000111011000;
rgb[3886] = 24'b111011101111000011101011;
rgb[3887] = 24'b111111111111111111111111;
rgb[3888] = 24'b000000000000000000000000;
rgb[3889] = 24'b000100010001010000001101;
rgb[3890] = 24'b001000100010100000011011;
rgb[3891] = 24'b001101000011110100101000;
rgb[3892] = 24'b010001010101000100110110;
rgb[3893] = 24'b010101110110010101000100;
rgb[3894] = 24'b011010000111101001010001;
rgb[3895] = 24'b011110101000111001011111;
rgb[3896] = 24'b100010111001111101110000;
rgb[3897] = 24'b100110111010110110000100;
rgb[3898] = 24'b101011001011101110011000;
rgb[3899] = 24'b101111001100100010101101;
rgb[3900] = 24'b110011011101011011000001;
rgb[3901] = 24'b110111011110001111010110;
rgb[3902] = 24'b111011101111000111101010;
rgb[3903] = 24'b111111111111111111111111;
rgb[3904] = 24'b000000000000000000000000;
rgb[3905] = 24'b000100010001010100001100;
rgb[3906] = 24'b001000110010101100011000;
rgb[3907] = 24'b001101000100000000100101;
rgb[3908] = 24'b010001100101011000110001;
rgb[3909] = 24'b010110000110101100111110;
rgb[3910] = 24'b011010011000000101001010;
rgb[3911] = 24'b011110111001011001010111;
rgb[3912] = 24'b100011001010011101101000;
rgb[3913] = 24'b100111001011010001111101;
rgb[3914] = 24'b101011011100000010010011;
rgb[3915] = 24'b101111011100110110101000;
rgb[3916] = 24'b110011011101100110111110;
rgb[3917] = 24'b110111101110011011010011;
rgb[3918] = 24'b111011101111001011101001;
rgb[3919] = 24'b111111111111111111111111;
rgb[3920] = 24'b000000000000000000000000;
rgb[3921] = 24'b000100010001011000001011;
rgb[3922] = 24'b001000110010110100010110;
rgb[3923] = 24'b001101010100010000100010;
rgb[3924] = 24'b010001110101101000101101;
rgb[3925] = 24'b010110010111000100111000;
rgb[3926] = 24'b011010101000100001000100;
rgb[3927] = 24'b011111001001111001001111;
rgb[3928] = 24'b100011011010111101100000;
rgb[3929] = 24'b100111011011101101110110;
rgb[3930] = 24'b101011101100011010001101;
rgb[3931] = 24'b101111101101000110100100;
rgb[3932] = 24'b110011101101110110111011;
rgb[3933] = 24'b110111101110100011010001;
rgb[3934] = 24'b111011101111001111101000;
rgb[3935] = 24'b111111111111111111111111;
rgb[3936] = 24'b000000000000000000000000;
rgb[3937] = 24'b000100010001011100001010;
rgb[3938] = 24'b001000110010111100010100;
rgb[3939] = 24'b001101010100011100011110;
rgb[3940] = 24'b010001110101111100101000;
rgb[3941] = 24'b010110010111011000110011;
rgb[3942] = 24'b011010111000111000111101;
rgb[3943] = 24'b011111011010011001000111;
rgb[3944] = 24'b100011101011011101011000;
rgb[3945] = 24'b100111101100000101110000;
rgb[3946] = 24'b101011101100110010000111;
rgb[3947] = 24'b101111101101011010011111;
rgb[3948] = 24'b110011101110000010110111;
rgb[3949] = 24'b110111101110101011001111;
rgb[3950] = 24'b111011101111010011100111;
rgb[3951] = 24'b111111101111111011111111;
rgb[3952] = 24'b000000000000000000000000;
rgb[3953] = 24'b000100100001100000001001;
rgb[3954] = 24'b001001000011000100010010;
rgb[3955] = 24'b001101100100101000011011;
rgb[3956] = 24'b010010000110001100100100;
rgb[3957] = 24'b010110100111110000101101;
rgb[3958] = 24'b011011001001010100110110;
rgb[3959] = 24'b011111101010111000111111;
rgb[3960] = 24'b100011111011111101010000;
rgb[3961] = 24'b100111111100100001101001;
rgb[3962] = 24'b101011111101000110000010;
rgb[3963] = 24'b101111111101101010011011;
rgb[3964] = 24'b110011111110001110110100;
rgb[3965] = 24'b110111111110110011001101;
rgb[3966] = 24'b111011111111010111100110;
rgb[3967] = 24'b111111111111111111111111;
rgb[3968] = 24'b000000000000000000000000;
rgb[3969] = 24'b000100100001101000000111;
rgb[3970] = 24'b001001000011010000001111;
rgb[3971] = 24'b001101100100111000010111;
rgb[3972] = 24'b010010010110100000011111;
rgb[3973] = 24'b010110111000001000100111;
rgb[3974] = 24'b011011011001110000101111;
rgb[3975] = 24'b100000001011011000110111;
rgb[3976] = 24'b100100011100011101001000;
rgb[3977] = 24'b101000001100111101100010;
rgb[3978] = 24'b101100001101011101111100;
rgb[3979] = 24'b110000001101111110010110;
rgb[3980] = 24'b110011111110011110110000;
rgb[3981] = 24'b110111111110111111001010;
rgb[3982] = 24'b111011111111011111100100;
rgb[3983] = 24'b111111101111111011111111;
rgb[3984] = 24'b000000000000000000000000;
rgb[3985] = 24'b000100100001101100000110;
rgb[3986] = 24'b001001000011011000001101;
rgb[3987] = 24'b001101110101000100010100;
rgb[3988] = 24'b010010010110110000011011;
rgb[3989] = 24'b010111001000100000100001;
rgb[3990] = 24'b011011101010001100101000;
rgb[3991] = 24'b100000011011111000101111;
rgb[3992] = 24'b100100101100111101000000;
rgb[3993] = 24'b101000011101011001011011;
rgb[3994] = 24'b101100011101110101110110;
rgb[3995] = 24'b110000001110001110010010;
rgb[3996] = 24'b110100001110101010101101;
rgb[3997] = 24'b110111111111000111001000;
rgb[3998] = 24'b111011111111100011100011;
rgb[3999] = 24'b111111111111111111111111;
rgb[4000] = 24'b000000000000000000000000;
rgb[4001] = 24'b000100100001110000000101;
rgb[4002] = 24'b001001010011100000001011;
rgb[4003] = 24'b001101110101010100010001;
rgb[4004] = 24'b010010100111000100010110;
rgb[4005] = 24'b010111011000110100011100;
rgb[4006] = 24'b011011111010101000100010;
rgb[4007] = 24'b100000101100011000100111;
rgb[4008] = 24'b100100111101011100111000;
rgb[4009] = 24'b101000101101110101010100;
rgb[4010] = 24'b101100101110001001110001;
rgb[4011] = 24'b110000011110100010001101;
rgb[4012] = 24'b110100001110111010101010;
rgb[4013] = 24'b111000001111001111000110;
rgb[4014] = 24'b111011111111100111100010;
rgb[4015] = 24'b111111101111111011111111;
rgb[4016] = 24'b000000000000000000000000;
rgb[4017] = 24'b000100100001110100000100;
rgb[4018] = 24'b001001010011101000001001;
rgb[4019] = 24'b001110000101100000001101;
rgb[4020] = 24'b010010110111010100010010;
rgb[4021] = 24'b010111011001001100010110;
rgb[4022] = 24'b011100001011000000011011;
rgb[4023] = 24'b100000111100111000011111;
rgb[4024] = 24'b100101001101111100110000;
rgb[4025] = 24'b101000111110001101001110;
rgb[4026] = 24'b101100101110100001101011;
rgb[4027] = 24'b110000101110110010001001;
rgb[4028] = 24'b110100011111000110100110;
rgb[4029] = 24'b111000001111010111000100;
rgb[4030] = 24'b111011111111101011100001;
rgb[4031] = 24'b111111111111111111111111;
rgb[4032] = 24'b000000000000000000000000;
rgb[4033] = 24'b000100100001111000000011;
rgb[4034] = 24'b001001010011110100000110;
rgb[4035] = 24'b001110000101101100001010;
rgb[4036] = 24'b010010110111101000001101;
rgb[4037] = 24'b010111101001100100010000;
rgb[4038] = 24'b011100011011011100010100;
rgb[4039] = 24'b100001001101011000010111;
rgb[4040] = 24'b100101011110011100101000;
rgb[4041] = 24'b101001001110101001000111;
rgb[4042] = 24'b101100111110111001100101;
rgb[4043] = 24'b110000101111000110000100;
rgb[4044] = 24'b110100011111010010100011;
rgb[4045] = 24'b111000001111100011000001;
rgb[4046] = 24'b111011111111101111100000;
rgb[4047] = 24'b111111111111111111111111;
rgb[4048] = 24'b000000000000000000000000;
rgb[4049] = 24'b000100110001111100000010;
rgb[4050] = 24'b001001100011111100000100;
rgb[4051] = 24'b001110010101111100000110;
rgb[4052] = 24'b010011000111111000001001;
rgb[4053] = 24'b010111111001111000001011;
rgb[4054] = 24'b011100101011111000001101;
rgb[4055] = 24'b100001011101111000001111;
rgb[4056] = 24'b100101101110111100100000;
rgb[4057] = 24'b101001011111000101000000;
rgb[4058] = 24'b101101001111001101100000;
rgb[4059] = 24'b110000111111010110000000;
rgb[4060] = 24'b110100101111100010011111;
rgb[4061] = 24'b111000011111101010111111;
rgb[4062] = 24'b111100001111110011011111;
rgb[4063] = 24'b111111111111111111111111;
rgb[4064] = 24'b000000000000000000000000;
rgb[4065] = 24'b000100110010000000000001;
rgb[4066] = 24'b001001100100000100000010;
rgb[4067] = 24'b001110010110001000000011;
rgb[4068] = 24'b010011011000001100000100;
rgb[4069] = 24'b011000001010010000000101;
rgb[4070] = 24'b011100111100010100000110;
rgb[4071] = 24'b100001101110011000000111;
rgb[4072] = 24'b100101111111011100011000;
rgb[4073] = 24'b101001101111100000111001;
rgb[4074] = 24'b101101011111100101011010;
rgb[4075] = 24'b110001001111101001111011;
rgb[4076] = 24'b110100101111101110011100;
rgb[4077] = 24'b111000011111110010111101;
rgb[4078] = 24'b111100001111110111011110;
rgb[4079] = 24'b111111111111111111111111;
rgb[4080] = 24'b000000000000000000000000;
rgb[4081] = 24'b000100110010001000000000;
rgb[4082] = 24'b001001100100010000000000;
rgb[4083] = 24'b001110100110011000000000;
rgb[4084] = 24'b010011011000100000000000;
rgb[4085] = 24'b011000011010101000000000;
rgb[4086] = 24'b011101001100110000000000;
rgb[4087] = 24'b100010001110111000000000;
rgb[4088] = 24'b100110011111111000010001;
rgb[4089] = 24'b101001111111111100110010;
rgb[4090] = 24'b101101101111111001010101;
rgb[4091] = 24'b110001001111111101110110;
rgb[4092] = 24'b110100111111111110011001;
rgb[4093] = 24'b111000011111111110111011;
rgb[4094] = 24'b111100001111111111011101;
rgb[4095] = 24'b111111111111111111111111;
rgb[4096] = 24'b000000000000000000000000;
rgb[4097] = 24'b000100010001000100010001;
rgb[4098] = 24'b001000100010001000100010;
rgb[4099] = 24'b001100110011001100110011;
rgb[4100] = 24'b010001000100010001000100;
rgb[4101] = 24'b010101010101010101010101;
rgb[4102] = 24'b011001100110011001100110;
rgb[4103] = 24'b011101110111011101110111;
rgb[4104] = 24'b100010001000100010001000;
rgb[4105] = 24'b100110011001100110011001;
rgb[4106] = 24'b101010101010101010101010;
rgb[4107] = 24'b101110111011101110111011;
rgb[4108] = 24'b110011001100110011001100;
rgb[4109] = 24'b110111011101110111011101;
rgb[4110] = 24'b111011101110111011101110;
rgb[4111] = 24'b111111111111111111111111;
rgb[4112] = 24'b000000000000000000000000;
rgb[4113] = 24'b000100000001001000001111;
rgb[4114] = 24'b001000010010010000011111;
rgb[4115] = 24'b001100100011011000101111;
rgb[4116] = 24'b010000110100100000111111;
rgb[4117] = 24'b010101000101101001001111;
rgb[4118] = 24'b011001010110110001011111;
rgb[4119] = 24'b011101100111111001101111;
rgb[4120] = 24'b100001111000111110000000;
rgb[4121] = 24'b100110001001111110010010;
rgb[4122] = 24'b101010011010111110100100;
rgb[4123] = 24'b101110101011111110110110;
rgb[4124] = 24'b110010111100111111001000;
rgb[4125] = 24'b110111001101111111011010;
rgb[4126] = 24'b111011011110111111101100;
rgb[4127] = 24'b111111111111111111111111;
rgb[4128] = 24'b000000000000000000000000;
rgb[4129] = 24'b000100000001001100001110;
rgb[4130] = 24'b001000010010011000011101;
rgb[4131] = 24'b001100100011100100101100;
rgb[4132] = 24'b010000110100110100111010;
rgb[4133] = 24'b010101000110000001001001;
rgb[4134] = 24'b011001010111001101011000;
rgb[4135] = 24'b011101101000011001100111;
rgb[4136] = 24'b100001111001011101111000;
rgb[4137] = 24'b100110001010011010001011;
rgb[4138] = 24'b101010011011010110011110;
rgb[4139] = 24'b101110101100010010110001;
rgb[4140] = 24'b110010111101001011000101;
rgb[4141] = 24'b110111001110000111011000;
rgb[4142] = 24'b111011011111000011101011;
rgb[4143] = 24'b111111111111111111111111;
rgb[4144] = 24'b000000000000000000000000;
rgb[4145] = 24'b000100000001010000001101;
rgb[4146] = 24'b001000010010100000011011;
rgb[4147] = 24'b001100100011110100101000;
rgb[4148] = 24'b010000110101000100110110;
rgb[4149] = 24'b010101000110010101000100;
rgb[4150] = 24'b011001010111101001010001;
rgb[4151] = 24'b011101011000111001011111;
rgb[4152] = 24'b100001101001111101110000;
rgb[4153] = 24'b100110001010110110000100;
rgb[4154] = 24'b101010011011101110011000;
rgb[4155] = 24'b101110101100100010101101;
rgb[4156] = 24'b110010111101011011000001;
rgb[4157] = 24'b110111001110001111010110;
rgb[4158] = 24'b111011011111000111101010;
rgb[4159] = 24'b111111111111111111111111;
rgb[4160] = 24'b000000000000000000000000;
rgb[4161] = 24'b000100000001010100001100;
rgb[4162] = 24'b001000010010101100011000;
rgb[4163] = 24'b001100100100000000100101;
rgb[4164] = 24'b010000110101011000110001;
rgb[4165] = 24'b010100110110101100111110;
rgb[4166] = 24'b011001001000000101001010;
rgb[4167] = 24'b011101011001011001010111;
rgb[4168] = 24'b100001101010011101101000;
rgb[4169] = 24'b100101111011010001111101;
rgb[4170] = 24'b101010001100000010010011;
rgb[4171] = 24'b101110101100110110101000;
rgb[4172] = 24'b110010111101100110111110;
rgb[4173] = 24'b110111001110011011010011;
rgb[4174] = 24'b111011011111001011101001;
rgb[4175] = 24'b111111111111111111111111;
rgb[4176] = 24'b000000000000000000000000;
rgb[4177] = 24'b000100000001011000001011;
rgb[4178] = 24'b001000010010110100010110;
rgb[4179] = 24'b001100100100010000100010;
rgb[4180] = 24'b010000100101101000101101;
rgb[4181] = 24'b010100110111000100111000;
rgb[4182] = 24'b011001001000100001000100;
rgb[4183] = 24'b011101011001111001001111;
rgb[4184] = 24'b100001101010111101100000;
rgb[4185] = 24'b100101111011101101110110;
rgb[4186] = 24'b101010001100011010001101;
rgb[4187] = 24'b101110011101000110100100;
rgb[4188] = 24'b110010111101110110111011;
rgb[4189] = 24'b110111001110100011010001;
rgb[4190] = 24'b111011011111001111101000;
rgb[4191] = 24'b111111111111111111111111;
rgb[4192] = 24'b000000000000000000000000;
rgb[4193] = 24'b000100000001011100001010;
rgb[4194] = 24'b001000010010111100010100;
rgb[4195] = 24'b001100100100011100011110;
rgb[4196] = 24'b010000100101111100101000;
rgb[4197] = 24'b010100110111011000110011;
rgb[4198] = 24'b011001001000111000111101;
rgb[4199] = 24'b011101001010011001000111;
rgb[4200] = 24'b100001011011011101011000;
rgb[4201] = 24'b100101111100000101110000;
rgb[4202] = 24'b101010001100110010000111;
rgb[4203] = 24'b101110011101011010011111;
rgb[4204] = 24'b110010111110000010110111;
rgb[4205] = 24'b110111001110101011001111;
rgb[4206] = 24'b111011011111010011100111;
rgb[4207] = 24'b111111111111111011111111;
rgb[4208] = 24'b000000000000000000000000;
rgb[4209] = 24'b000100000001100000001001;
rgb[4210] = 24'b001000010011000100010010;
rgb[4211] = 24'b001100010100101000011011;
rgb[4212] = 24'b010000100110001100100100;
rgb[4213] = 24'b010100110111110000101101;
rgb[4214] = 24'b011000111001010100110110;
rgb[4215] = 24'b011101001010111000111111;
rgb[4216] = 24'b100001011011111101010000;
rgb[4217] = 24'b100101101100100001101001;
rgb[4218] = 24'b101010001101000110000010;
rgb[4219] = 24'b101110011101101010011011;
rgb[4220] = 24'b110010101110001110110100;
rgb[4221] = 24'b110111001110110011001101;
rgb[4222] = 24'b111011011111010111100110;
rgb[4223] = 24'b111111111111111111111111;
rgb[4224] = 24'b000000000000000000000000;
rgb[4225] = 24'b000100000001101000000111;
rgb[4226] = 24'b001000010011010000001111;
rgb[4227] = 24'b001100010100111000010111;
rgb[4228] = 24'b010000100110100000011111;
rgb[4229] = 24'b010100101000001000100111;
rgb[4230] = 24'b011000111001110000101111;
rgb[4231] = 24'b011100111011011000110111;
rgb[4232] = 24'b100001001100011101001000;
rgb[4233] = 24'b100101101100111101100010;
rgb[4234] = 24'b101001111101011101111100;
rgb[4235] = 24'b101110011101111110010110;
rgb[4236] = 24'b110010101110011110110000;
rgb[4237] = 24'b110111001110111111001010;
rgb[4238] = 24'b111011011111011111100100;
rgb[4239] = 24'b111111111111111011111111;
rgb[4240] = 24'b000000000000000000000000;
rgb[4241] = 24'b000100000001101100000110;
rgb[4242] = 24'b001000010011011000001101;
rgb[4243] = 24'b001100010101000100010100;
rgb[4244] = 24'b010000100110110000011011;
rgb[4245] = 24'b010100101000100000100001;
rgb[4246] = 24'b011000111010001100101000;
rgb[4247] = 24'b011100111011111000101111;
rgb[4248] = 24'b100001001100111101000000;
rgb[4249] = 24'b100101101101011001011011;
rgb[4250] = 24'b101001111101110101110110;
rgb[4251] = 24'b101110011110001110010010;
rgb[4252] = 24'b110010101110101010101101;
rgb[4253] = 24'b110111001111000111001000;
rgb[4254] = 24'b111011011111100011100011;
rgb[4255] = 24'b111111111111111111111111;
rgb[4256] = 24'b000000000000000000000000;
rgb[4257] = 24'b000100000001110000000101;
rgb[4258] = 24'b001000000011100000001011;
rgb[4259] = 24'b001100010101010100010001;
rgb[4260] = 24'b010000010111000100010110;
rgb[4261] = 24'b010100101000110100011100;
rgb[4262] = 24'b011000101010101000100010;
rgb[4263] = 24'b011100111100011000100111;
rgb[4264] = 24'b100001001101011100111000;
rgb[4265] = 24'b100101011101110101010100;
rgb[4266] = 24'b101001111110001001110001;
rgb[4267] = 24'b101110001110100010001101;
rgb[4268] = 24'b110010101110111010101010;
rgb[4269] = 24'b110110111111001111000110;
rgb[4270] = 24'b111011011111100111100010;
rgb[4271] = 24'b111111111111111011111111;
rgb[4272] = 24'b000000000000000000000000;
rgb[4273] = 24'b000100000001110100000100;
rgb[4274] = 24'b001000000011101000001001;
rgb[4275] = 24'b001100010101100000001101;
rgb[4276] = 24'b010000010111010100010010;
rgb[4277] = 24'b010100101001001100010110;
rgb[4278] = 24'b011000101011000000011011;
rgb[4279] = 24'b011100101100111000011111;
rgb[4280] = 24'b100000111101111100110000;
rgb[4281] = 24'b100101011110001101001110;
rgb[4282] = 24'b101001111110100001101011;
rgb[4283] = 24'b101110001110110010001001;
rgb[4284] = 24'b110010101111000110100110;
rgb[4285] = 24'b110110111111010111000100;
rgb[4286] = 24'b111011011111101011100001;
rgb[4287] = 24'b111111111111111111111111;
rgb[4288] = 24'b000000000000000000000000;
rgb[4289] = 24'b000100000001111000000011;
rgb[4290] = 24'b001000000011110100000110;
rgb[4291] = 24'b001100010101101100001010;
rgb[4292] = 24'b010000010111101000001101;
rgb[4293] = 24'b010100011001100100010000;
rgb[4294] = 24'b011000101011011100010100;
rgb[4295] = 24'b011100101101011000010111;
rgb[4296] = 24'b100000111110011100101000;
rgb[4297] = 24'b100101011110101001000111;
rgb[4298] = 24'b101001101110111001100101;
rgb[4299] = 24'b101110001111000110000100;
rgb[4300] = 24'b110010101111010010100011;
rgb[4301] = 24'b110110111111100011000001;
rgb[4302] = 24'b111011011111101111100000;
rgb[4303] = 24'b111111111111111111111111;
rgb[4304] = 24'b000000000000000000000000;
rgb[4305] = 24'b000100000001111100000010;
rgb[4306] = 24'b001000000011111100000100;
rgb[4307] = 24'b001100000101111100000110;
rgb[4308] = 24'b010000010111111000001001;
rgb[4309] = 24'b010100011001111000001011;
rgb[4310] = 24'b011000011011111000001101;
rgb[4311] = 24'b011100101101111000001111;
rgb[4312] = 24'b100000111110111100100000;
rgb[4313] = 24'b100101001111000101000000;
rgb[4314] = 24'b101001101111001101100000;
rgb[4315] = 24'b101110001111010110000000;
rgb[4316] = 24'b110010011111100010011111;
rgb[4317] = 24'b110110111111101010111111;
rgb[4318] = 24'b111011011111110011011111;
rgb[4319] = 24'b111111111111111111111111;
rgb[4320] = 24'b000000000000000000000000;
rgb[4321] = 24'b000100000010000000000001;
rgb[4322] = 24'b001000000100000100000010;
rgb[4323] = 24'b001100000110001000000011;
rgb[4324] = 24'b010000001000001100000100;
rgb[4325] = 24'b010100011010010000000101;
rgb[4326] = 24'b011000011100010100000110;
rgb[4327] = 24'b011100011110011000000111;
rgb[4328] = 24'b100000101111011100011000;
rgb[4329] = 24'b100101001111100000111001;
rgb[4330] = 24'b101001101111100101011010;
rgb[4331] = 24'b101101111111101001111011;
rgb[4332] = 24'b110010011111101110011100;
rgb[4333] = 24'b110110111111110010111101;
rgb[4334] = 24'b111011011111110111011110;
rgb[4335] = 24'b111111111111111111111111;
rgb[4336] = 24'b000000000000000000000000;
rgb[4337] = 24'b000100000010001000000000;
rgb[4338] = 24'b001000000100010000000000;
rgb[4339] = 24'b001100000110011000000000;
rgb[4340] = 24'b010000001000100000000000;
rgb[4341] = 24'b010100001010101000000000;
rgb[4342] = 24'b011000011100110000000000;
rgb[4343] = 24'b011100011110111000000000;
rgb[4344] = 24'b100000101111111000010001;
rgb[4345] = 24'b100101001111111100110010;
rgb[4346] = 24'b101001011111111001010101;
rgb[4347] = 24'b101101111111111101110110;
rgb[4348] = 24'b110010011111111110011001;
rgb[4349] = 24'b110110111111111110111011;
rgb[4350] = 24'b111011011111111111011101;
rgb[4351] = 24'b111111111111111111111111;
rgb[4352] = 24'b000000000000000000000000;
rgb[4353] = 24'b000100010001000100010001;
rgb[4354] = 24'b001000100010001000100010;
rgb[4355] = 24'b001100110011001100110011;
rgb[4356] = 24'b010001000100010001000100;
rgb[4357] = 24'b010101010101010101010101;
rgb[4358] = 24'b011001100110011001100110;
rgb[4359] = 24'b011101110111011101110111;
rgb[4360] = 24'b100010001000100010001000;
rgb[4361] = 24'b100110011001100110011001;
rgb[4362] = 24'b101010101010101010101010;
rgb[4363] = 24'b101110111011101110111011;
rgb[4364] = 24'b110011001100110011001100;
rgb[4365] = 24'b110111011101110111011101;
rgb[4366] = 24'b111011101110111011101110;
rgb[4367] = 24'b111111111111111111111111;
rgb[4368] = 24'b000000000000000000000000;
rgb[4369] = 24'b000100000001001000001111;
rgb[4370] = 24'b001000010010010000011111;
rgb[4371] = 24'b001100100011011000101111;
rgb[4372] = 24'b010000100100100000111111;
rgb[4373] = 24'b010100110101101001001111;
rgb[4374] = 24'b011001000110110001011111;
rgb[4375] = 24'b011101010111111001101111;
rgb[4376] = 24'b100001101000111110000000;
rgb[4377] = 24'b100101111001111110010010;
rgb[4378] = 24'b101010001010111110100100;
rgb[4379] = 24'b101110011011111110110110;
rgb[4380] = 24'b110010111100111111001000;
rgb[4381] = 24'b110111001101111111011010;
rgb[4382] = 24'b111011011110111111101100;
rgb[4383] = 24'b111111111111111111111111;
rgb[4384] = 24'b000000000000000000000000;
rgb[4385] = 24'b000100000001001100001110;
rgb[4386] = 24'b001000000010011000011101;
rgb[4387] = 24'b001100010011100100101100;
rgb[4388] = 24'b010000010100110100111010;
rgb[4389] = 24'b010100100110000001001001;
rgb[4390] = 24'b011000100111001101011000;
rgb[4391] = 24'b011100111000011001100111;
rgb[4392] = 24'b100001001001011101111000;
rgb[4393] = 24'b100101011010011010001011;
rgb[4394] = 24'b101001111011010110011110;
rgb[4395] = 24'b101110001100010010110001;
rgb[4396] = 24'b110010101101001011000101;
rgb[4397] = 24'b110110111110000111011000;
rgb[4398] = 24'b111011011111000011101011;
rgb[4399] = 24'b111111111111111111111111;
rgb[4400] = 24'b000000000000000000000000;
rgb[4401] = 24'b000100000001010000001101;
rgb[4402] = 24'b001000000010100000011011;
rgb[4403] = 24'b001100000011110100101000;
rgb[4404] = 24'b010000000101000100110110;
rgb[4405] = 24'b010100000110010101000100;
rgb[4406] = 24'b011000010111101001010001;
rgb[4407] = 24'b011100011000111001011111;
rgb[4408] = 24'b100000101001111101110000;
rgb[4409] = 24'b100101001010110110000100;
rgb[4410] = 24'b101001011011101110011000;
rgb[4411] = 24'b101101111100100010101101;
rgb[4412] = 24'b110010011101011011000001;
rgb[4413] = 24'b110110111110001111010110;
rgb[4414] = 24'b111011011111000111101010;
rgb[4415] = 24'b111111111111111111111111;
rgb[4416] = 24'b000000000000000000000000;
rgb[4417] = 24'b000011110001010100001100;
rgb[4418] = 24'b000111110010101100011000;
rgb[4419] = 24'b001011110100000000100101;
rgb[4420] = 24'b001111110101011000110001;
rgb[4421] = 24'b010011110110101100111110;
rgb[4422] = 24'b010111111000000101001010;
rgb[4423] = 24'b011011111001011001010111;
rgb[4424] = 24'b100000001010011101101000;
rgb[4425] = 24'b100100101011010001111101;
rgb[4426] = 24'b101001001100000010010011;
rgb[4427] = 24'b101101101100110110101000;
rgb[4428] = 24'b110010001101100110111110;
rgb[4429] = 24'b110110101110011011010011;
rgb[4430] = 24'b111011001111001011101001;
rgb[4431] = 24'b111111111111111111111111;
rgb[4432] = 24'b000000000000000000000000;
rgb[4433] = 24'b000011110001011000001011;
rgb[4434] = 24'b000111110010110100010110;
rgb[4435] = 24'b001011100100010000100010;
rgb[4436] = 24'b001111100101101000101101;
rgb[4437] = 24'b010011100111000100111000;
rgb[4438] = 24'b010111011000100001000100;
rgb[4439] = 24'b011011011001111001001111;
rgb[4440] = 24'b011111101010111101100000;
rgb[4441] = 24'b100100001011101101110110;
rgb[4442] = 24'b101000111100011010001101;
rgb[4443] = 24'b101101011101000110100100;
rgb[4444] = 24'b110001111101110110111011;
rgb[4445] = 24'b110110101110100011010001;
rgb[4446] = 24'b111011001111001111101000;
rgb[4447] = 24'b111111111111111111111111;
rgb[4448] = 24'b000000000000000000000000;
rgb[4449] = 24'b000011110001011100001010;
rgb[4450] = 24'b000111100010111100010100;
rgb[4451] = 24'b001011100100011100011110;
rgb[4452] = 24'b001111010101111100101000;
rgb[4453] = 24'b010011000111011000110011;
rgb[4454] = 24'b010111001000111000111101;
rgb[4455] = 24'b011010111010011001000111;
rgb[4456] = 24'b011111001011011101011000;
rgb[4457] = 24'b100011111100000101110000;
rgb[4458] = 24'b101000011100110010000111;
rgb[4459] = 24'b101101001101011010011111;
rgb[4460] = 24'b110001111110000010110111;
rgb[4461] = 24'b110110011110101011001111;
rgb[4462] = 24'b111011001111010011100111;
rgb[4463] = 24'b111111111111111011111111;
rgb[4464] = 24'b000000000000000000000000;
rgb[4465] = 24'b000011110001100000001001;
rgb[4466] = 24'b000111100011000100010010;
rgb[4467] = 24'b001011010100101000011011;
rgb[4468] = 24'b001111000110001100100100;
rgb[4469] = 24'b010010110111110000101101;
rgb[4470] = 24'b010110101001010100110110;
rgb[4471] = 24'b011010011010111000111111;
rgb[4472] = 24'b011110101011111101010000;
rgb[4473] = 24'b100011011100100001101001;
rgb[4474] = 24'b101000001101000110000010;
rgb[4475] = 24'b101100111101101010011011;
rgb[4476] = 24'b110001101110001110110100;
rgb[4477] = 24'b110110011110110011001101;
rgb[4478] = 24'b111011001111010111100110;
rgb[4479] = 24'b111111111111111111111111;
rgb[4480] = 24'b000000000000000000000000;
rgb[4481] = 24'b000011100001101000000111;
rgb[4482] = 24'b000111010011010000001111;
rgb[4483] = 24'b001011000100111000010111;
rgb[4484] = 24'b001110110110100000011111;
rgb[4485] = 24'b010010101000001000100111;
rgb[4486] = 24'b010110011001110000101111;
rgb[4487] = 24'b011001111011011000110111;
rgb[4488] = 24'b011110001100011101001000;
rgb[4489] = 24'b100011001100111101100010;
rgb[4490] = 24'b100111111101011101111100;
rgb[4491] = 24'b101100101101111110010110;
rgb[4492] = 24'b110001011110011110110000;
rgb[4493] = 24'b110110001110111111001010;
rgb[4494] = 24'b111010111111011111100100;
rgb[4495] = 24'b111111111111111011111111;
rgb[4496] = 24'b000000000000000000000000;
rgb[4497] = 24'b000011100001101100000110;
rgb[4498] = 24'b000111010011011000001101;
rgb[4499] = 24'b001010110101000100010100;
rgb[4500] = 24'b001110100110110000011011;
rgb[4501] = 24'b010010001000100000100001;
rgb[4502] = 24'b010101111010001100101000;
rgb[4503] = 24'b011001011011111000101111;
rgb[4504] = 24'b011101111100111101000000;
rgb[4505] = 24'b100010101101011001011011;
rgb[4506] = 24'b100111011101110101110110;
rgb[4507] = 24'b101100011110001110010010;
rgb[4508] = 24'b110001001110101010101101;
rgb[4509] = 24'b110110001111000111001000;
rgb[4510] = 24'b111010111111100011100011;
rgb[4511] = 24'b111111111111111111111111;
rgb[4512] = 24'b000000000000000000000000;
rgb[4513] = 24'b000011100001110000000101;
rgb[4514] = 24'b000111000011100000001011;
rgb[4515] = 24'b001010100101010100010001;
rgb[4516] = 24'b001110010111000100010110;
rgb[4517] = 24'b010001111000110100011100;
rgb[4518] = 24'b010101011010101000100010;
rgb[4519] = 24'b011001001100011000100111;
rgb[4520] = 24'b011101011101011100111000;
rgb[4521] = 24'b100010001101110101010100;
rgb[4522] = 24'b100111001110001001110001;
rgb[4523] = 24'b101100001110100010001101;
rgb[4524] = 24'b110000111110111010101010;
rgb[4525] = 24'b110101111111001111000110;
rgb[4526] = 24'b111010111111100111100010;
rgb[4527] = 24'b111111111111111011111111;
rgb[4528] = 24'b000000000000000000000000;
rgb[4529] = 24'b000011100001110100000100;
rgb[4530] = 24'b000111000011101000001001;
rgb[4531] = 24'b001010100101100000001101;
rgb[4532] = 24'b001110000111010100010010;
rgb[4533] = 24'b010001101001001100010110;
rgb[4534] = 24'b010101001011000000011011;
rgb[4535] = 24'b011000101100111000011111;
rgb[4536] = 24'b011100111101111100110000;
rgb[4537] = 24'b100001111110001101001110;
rgb[4538] = 24'b100110111110100001101011;
rgb[4539] = 24'b101011111110110010001001;
rgb[4540] = 24'b110000111111000110100110;
rgb[4541] = 24'b110101111111010111000100;
rgb[4542] = 24'b111010111111101011100001;
rgb[4543] = 24'b111111111111111111111111;
rgb[4544] = 24'b000000000000000000000000;
rgb[4545] = 24'b000011010001111000000011;
rgb[4546] = 24'b000110110011110100000110;
rgb[4547] = 24'b001010010101101100001010;
rgb[4548] = 24'b001101110111101000001101;
rgb[4549] = 24'b010001001001100100010000;
rgb[4550] = 24'b010100101011011100010100;
rgb[4551] = 24'b011000001101011000010111;
rgb[4552] = 24'b011100011110011100101000;
rgb[4553] = 24'b100001011110101001000111;
rgb[4554] = 24'b100110011110111001100101;
rgb[4555] = 24'b101011101111000110000100;
rgb[4556] = 24'b110000101111010010100011;
rgb[4557] = 24'b110101101111100011000001;
rgb[4558] = 24'b111010101111101111100000;
rgb[4559] = 24'b111111111111111111111111;
rgb[4560] = 24'b000000000000000000000000;
rgb[4561] = 24'b000011010001111100000010;
rgb[4562] = 24'b000110100011111100000100;
rgb[4563] = 24'b001010000101111100000110;
rgb[4564] = 24'b001101010111111000001001;
rgb[4565] = 24'b010000111001111000001011;
rgb[4566] = 24'b010100001011111000001101;
rgb[4567] = 24'b010111101101111000001111;
rgb[4568] = 24'b011011111110111100100000;
rgb[4569] = 24'b100000111111000101000000;
rgb[4570] = 24'b100110001111001101100000;
rgb[4571] = 24'b101011001111010110000000;
rgb[4572] = 24'b110000011111100010011111;
rgb[4573] = 24'b110101011111101010111111;
rgb[4574] = 24'b111010101111110011011111;
rgb[4575] = 24'b111111111111111111111111;
rgb[4576] = 24'b000000000000000000000000;
rgb[4577] = 24'b000011010010000000000001;
rgb[4578] = 24'b000110100100000100000010;
rgb[4579] = 24'b001001110110001000000011;
rgb[4580] = 24'b001101001000001100000100;
rgb[4581] = 24'b010000101010010000000101;
rgb[4582] = 24'b010011111100010100000110;
rgb[4583] = 24'b010111001110011000000111;
rgb[4584] = 24'b011011011111011100011000;
rgb[4585] = 24'b100000101111100000111001;
rgb[4586] = 24'b100101111111100101011010;
rgb[4587] = 24'b101010111111101001111011;
rgb[4588] = 24'b110000001111101110011100;
rgb[4589] = 24'b110101011111110010111101;
rgb[4590] = 24'b111010101111110111011110;
rgb[4591] = 24'b111111111111111111111111;
rgb[4592] = 24'b000000000000000000000000;
rgb[4593] = 24'b000011000010001000000000;
rgb[4594] = 24'b000110010100010000000000;
rgb[4595] = 24'b001001100110011000000000;
rgb[4596] = 24'b001100111000100000000000;
rgb[4597] = 24'b010000001010101000000000;
rgb[4598] = 24'b010011011100110000000000;
rgb[4599] = 24'b010110101110111000000000;
rgb[4600] = 24'b011010111111111000010001;
rgb[4601] = 24'b100000001111111100110010;
rgb[4602] = 24'b100101011111111001010101;
rgb[4603] = 24'b101010101111111101110110;
rgb[4604] = 24'b101111111111111110011001;
rgb[4605] = 24'b110101001111111110111011;
rgb[4606] = 24'b111010011111111111011101;
rgb[4607] = 24'b111111111111111111111111;
rgb[4608] = 24'b000000000000000000000000;
rgb[4609] = 24'b000100010001000100010001;
rgb[4610] = 24'b001000100010001000100010;
rgb[4611] = 24'b001100110011001100110011;
rgb[4612] = 24'b010001000100010001000100;
rgb[4613] = 24'b010101010101010101010101;
rgb[4614] = 24'b011001100110011001100110;
rgb[4615] = 24'b011101110111011101110111;
rgb[4616] = 24'b100010001000100010001000;
rgb[4617] = 24'b100110011001100110011001;
rgb[4618] = 24'b101010101010101010101010;
rgb[4619] = 24'b101110111011101110111011;
rgb[4620] = 24'b110011001100110011001100;
rgb[4621] = 24'b110111011101110111011101;
rgb[4622] = 24'b111011101110111011101110;
rgb[4623] = 24'b111111111111111111111111;
rgb[4624] = 24'b000000000000000000000000;
rgb[4625] = 24'b000100000001001000001111;
rgb[4626] = 24'b001000010010010000011111;
rgb[4627] = 24'b001100010011011000101111;
rgb[4628] = 24'b010000100100100000111111;
rgb[4629] = 24'b010100100101101001001111;
rgb[4630] = 24'b011000110110110001011111;
rgb[4631] = 24'b011100110111111001101111;
rgb[4632] = 24'b100001001000111110000000;
rgb[4633] = 24'b100101101001111110010010;
rgb[4634] = 24'b101001111010111110100100;
rgb[4635] = 24'b101110011011111110110110;
rgb[4636] = 24'b110010101100111111001000;
rgb[4637] = 24'b110111001101111111011010;
rgb[4638] = 24'b111011011110111111101100;
rgb[4639] = 24'b111111111111111111111111;
rgb[4640] = 24'b000000000000000000000000;
rgb[4641] = 24'b000100000001001100001110;
rgb[4642] = 24'b001000000010011000011101;
rgb[4643] = 24'b001100000011100100101100;
rgb[4644] = 24'b010000000100110100111010;
rgb[4645] = 24'b010100000110000001001001;
rgb[4646] = 24'b011000000111001101011000;
rgb[4647] = 24'b011100001000011001100111;
rgb[4648] = 24'b100000011001011101111000;
rgb[4649] = 24'b100100111010011010001011;
rgb[4650] = 24'b101001011011010110011110;
rgb[4651] = 24'b101101111100010010110001;
rgb[4652] = 24'b110010011101001011000101;
rgb[4653] = 24'b110110111110000111011000;
rgb[4654] = 24'b111011011111000011101011;
rgb[4655] = 24'b111111111111111111111111;
rgb[4656] = 24'b000000000000000000000000;
rgb[4657] = 24'b000011110001010000001101;
rgb[4658] = 24'b000111110010100000011011;
rgb[4659] = 24'b001011100011110100101000;
rgb[4660] = 24'b001111100101000100110110;
rgb[4661] = 24'b010011010110010101000100;
rgb[4662] = 24'b010111010111101001010001;
rgb[4663] = 24'b011011001000111001011111;
rgb[4664] = 24'b011111011001111101110000;
rgb[4665] = 24'b100100001010110110000100;
rgb[4666] = 24'b101000101011101110011000;
rgb[4667] = 24'b101101011100100010101101;
rgb[4668] = 24'b110001111101011011000001;
rgb[4669] = 24'b110110101110001111010110;
rgb[4670] = 24'b111011001111000111101010;
rgb[4671] = 24'b111111111111111111111111;
rgb[4672] = 24'b000000000000000000000000;
rgb[4673] = 24'b000011110001010100001100;
rgb[4674] = 24'b000111100010101100011000;
rgb[4675] = 24'b001011010100000000100101;
rgb[4676] = 24'b001111000101011000110001;
rgb[4677] = 24'b010010110110101100111110;
rgb[4678] = 24'b010110101000000101001010;
rgb[4679] = 24'b011010011001011001010111;
rgb[4680] = 24'b011110101010011101101000;
rgb[4681] = 24'b100011011011010001111101;
rgb[4682] = 24'b101000001100000010010011;
rgb[4683] = 24'b101100111100110110101000;
rgb[4684] = 24'b110001101101100110111110;
rgb[4685] = 24'b110110011110011011010011;
rgb[4686] = 24'b111011001111001011101001;
rgb[4687] = 24'b111111111111111111111111;
rgb[4688] = 24'b000000000000000000000000;
rgb[4689] = 24'b000011100001011000001011;
rgb[4690] = 24'b000111010010110100010110;
rgb[4691] = 24'b001010110100010000100010;
rgb[4692] = 24'b001110100101101000101101;
rgb[4693] = 24'b010010000111000100111000;
rgb[4694] = 24'b010101111000100001000100;
rgb[4695] = 24'b011001011001111001001111;
rgb[4696] = 24'b011101101010111101100000;
rgb[4697] = 24'b100010101011101101110110;
rgb[4698] = 24'b100111011100011010001101;
rgb[4699] = 24'b101100011101000110100100;
rgb[4700] = 24'b110001001101110110111011;
rgb[4701] = 24'b110110001110100011010001;
rgb[4702] = 24'b111010111111001111101000;
rgb[4703] = 24'b111111111111111111111111;
rgb[4704] = 24'b000000000000000000000000;
rgb[4705] = 24'b000011100001011100001010;
rgb[4706] = 24'b000111000010111100010100;
rgb[4707] = 24'b001010100100011100011110;
rgb[4708] = 24'b001110000101111100101000;
rgb[4709] = 24'b010001100111011000110011;
rgb[4710] = 24'b010101001000111000111101;
rgb[4711] = 24'b011000101010011001000111;
rgb[4712] = 24'b011100111011011101011000;
rgb[4713] = 24'b100001111100000101110000;
rgb[4714] = 24'b100110111100110010000111;
rgb[4715] = 24'b101011111101011010011111;
rgb[4716] = 24'b110000111110000010110111;
rgb[4717] = 24'b110101111110101011001111;
rgb[4718] = 24'b111010111111010011100111;
rgb[4719] = 24'b111111111111111011111111;
rgb[4720] = 24'b000000000000000000000000;
rgb[4721] = 24'b000011010001100000001001;
rgb[4722] = 24'b000110110011000100010010;
rgb[4723] = 24'b001010000100101000011011;
rgb[4724] = 24'b001101100110001100100100;
rgb[4725] = 24'b010000110111110000101101;
rgb[4726] = 24'b010100011001010100110110;
rgb[4727] = 24'b010111111010111000111111;
rgb[4728] = 24'b011100001011111101010000;
rgb[4729] = 24'b100001001100100001101001;
rgb[4730] = 24'b100110001101000110000010;
rgb[4731] = 24'b101011011101101010011011;
rgb[4732] = 24'b110000011110001110110100;
rgb[4733] = 24'b110101101110110011001101;
rgb[4734] = 24'b111010101111010111100110;
rgb[4735] = 24'b111111111111111111111111;
rgb[4736] = 24'b000000000000000000000000;
rgb[4737] = 24'b000011010001101000000111;
rgb[4738] = 24'b000110100011010000001111;
rgb[4739] = 24'b001001110100111000010111;
rgb[4740] = 24'b001101000110100000011111;
rgb[4741] = 24'b010000011000001000100111;
rgb[4742] = 24'b010011101001110000101111;
rgb[4743] = 24'b010110111011011000110111;
rgb[4744] = 24'b011011001100011101001000;
rgb[4745] = 24'b100000011100111101100010;
rgb[4746] = 24'b100101101101011101111100;
rgb[4747] = 24'b101010111101111110010110;
rgb[4748] = 24'b110000001110011110110000;
rgb[4749] = 24'b110101011110111111001010;
rgb[4750] = 24'b111010101111011111100100;
rgb[4751] = 24'b111111111111111011111111;
rgb[4752] = 24'b000000000000000000000000;
rgb[4753] = 24'b000011000001101100000110;
rgb[4754] = 24'b000110010011011000001101;
rgb[4755] = 24'b001001010101000100010100;
rgb[4756] = 24'b001100100110110000011011;
rgb[4757] = 24'b001111111000100000100001;
rgb[4758] = 24'b010010111010001100101000;
rgb[4759] = 24'b010110001011111000101111;
rgb[4760] = 24'b011010011100111101000000;
rgb[4761] = 24'b011111101101011001011011;
rgb[4762] = 24'b100101001101110101110110;
rgb[4763] = 24'b101010011110001110010010;
rgb[4764] = 24'b101111101110101010101101;
rgb[4765] = 24'b110101001111000111001000;
rgb[4766] = 24'b111010011111100011100011;
rgb[4767] = 24'b111111111111111111111111;
rgb[4768] = 24'b000000000000000000000000;
rgb[4769] = 24'b000011000001110000000101;
rgb[4770] = 24'b000110000011100000001011;
rgb[4771] = 24'b001001000101010100010001;
rgb[4772] = 24'b001100000111000100010110;
rgb[4773] = 24'b001111001000110100011100;
rgb[4774] = 24'b010010001010101000100010;
rgb[4775] = 24'b010101001100011000100111;
rgb[4776] = 24'b011001011101011100111000;
rgb[4777] = 24'b011110111101110101010100;
rgb[4778] = 24'b100100011110001001110001;
rgb[4779] = 24'b101001111110100010001101;
rgb[4780] = 24'b101111011110111010101010;
rgb[4781] = 24'b110100111111001111000110;
rgb[4782] = 24'b111010011111100111100010;
rgb[4783] = 24'b111111111111111011111111;
rgb[4784] = 24'b000000000000000000000000;
rgb[4785] = 24'b000010110001110100000100;
rgb[4786] = 24'b000101110011101000001001;
rgb[4787] = 24'b001000100101100000001101;
rgb[4788] = 24'b001011100111010100010010;
rgb[4789] = 24'b001110101001001100010110;
rgb[4790] = 24'b010001011011000000011011;
rgb[4791] = 24'b010100011100111000011111;
rgb[4792] = 24'b011000101101111100110000;
rgb[4793] = 24'b011110001110001101001110;
rgb[4794] = 24'b100011111110100001101011;
rgb[4795] = 24'b101001011110110010001001;
rgb[4796] = 24'b101110111111000110100110;
rgb[4797] = 24'b110100101111010111000100;
rgb[4798] = 24'b111010001111101011100001;
rgb[4799] = 24'b111111111111111111111111;
rgb[4800] = 24'b000000000000000000000000;
rgb[4801] = 24'b000010110001111000000011;
rgb[4802] = 24'b000101100011110100000110;
rgb[4803] = 24'b001000010101101100001010;
rgb[4804] = 24'b001011000111101000001101;
rgb[4805] = 24'b001101111001100100010000;
rgb[4806] = 24'b010000111011011100010100;
rgb[4807] = 24'b010011101101011000010111;
rgb[4808] = 24'b010111111110011100101000;
rgb[4809] = 24'b011101101110101001000111;
rgb[4810] = 24'b100011001110111001100101;
rgb[4811] = 24'b101000111111000110000100;
rgb[4812] = 24'b101110101111010010100011;
rgb[4813] = 24'b110100011111100011000001;
rgb[4814] = 24'b111010001111101111100000;
rgb[4815] = 24'b111111111111111111111111;
rgb[4816] = 24'b000000000000000000000000;
rgb[4817] = 24'b000010100001111100000010;
rgb[4818] = 24'b000101010011111100000100;
rgb[4819] = 24'b001000000101111100000110;
rgb[4820] = 24'b001010100111111000001001;
rgb[4821] = 24'b001101011001111000001011;
rgb[4822] = 24'b010000001011111000001101;
rgb[4823] = 24'b010010101101111000001111;
rgb[4824] = 24'b010110111110111100100000;
rgb[4825] = 24'b011100111111000101000000;
rgb[4826] = 24'b100010101111001101100000;
rgb[4827] = 24'b101000011111010110000000;
rgb[4828] = 24'b101110011111100010011111;
rgb[4829] = 24'b110100001111101010111111;
rgb[4830] = 24'b111001111111110011011111;
rgb[4831] = 24'b111111111111111111111111;
rgb[4832] = 24'b000000000000000000000000;
rgb[4833] = 24'b000010100010000000000001;
rgb[4834] = 24'b000101000100000100000010;
rgb[4835] = 24'b000111100110001000000011;
rgb[4836] = 24'b001010001000001100000100;
rgb[4837] = 24'b001100101010010000000101;
rgb[4838] = 24'b001111011100010100000110;
rgb[4839] = 24'b010001111110011000000111;
rgb[4840] = 24'b010110001111011100011000;
rgb[4841] = 24'b011100001111100000111001;
rgb[4842] = 24'b100001111111100101011010;
rgb[4843] = 24'b100111111111101001111011;
rgb[4844] = 24'b101101111111101110011100;
rgb[4845] = 24'b110011111111110010111101;
rgb[4846] = 24'b111001111111110111011110;
rgb[4847] = 24'b111111111111111111111111;
rgb[4848] = 24'b000000000000000000000000;
rgb[4849] = 24'b000010010010001000000000;
rgb[4850] = 24'b000100110100010000000000;
rgb[4851] = 24'b000111010110011000000000;
rgb[4852] = 24'b001001101000100000000000;
rgb[4853] = 24'b001100001010101000000000;
rgb[4854] = 24'b001110101100110000000000;
rgb[4855] = 24'b010000111110111000000000;
rgb[4856] = 24'b010101001111111000010001;
rgb[4857] = 24'b011011011111111100110010;
rgb[4858] = 24'b100001011111111001010101;
rgb[4859] = 24'b100111011111111101110110;
rgb[4860] = 24'b101101101111111110011001;
rgb[4861] = 24'b110011101111111110111011;
rgb[4862] = 24'b111001101111111111011101;
rgb[4863] = 24'b111111111111111111111111;
rgb[4864] = 24'b000000000000000000000000;
rgb[4865] = 24'b000100010001000100010001;
rgb[4866] = 24'b001000100010001000100010;
rgb[4867] = 24'b001100110011001100110011;
rgb[4868] = 24'b010001000100010001000100;
rgb[4869] = 24'b010101010101010101010101;
rgb[4870] = 24'b011001100110011001100110;
rgb[4871] = 24'b011101110111011101110111;
rgb[4872] = 24'b100010001000100010001000;
rgb[4873] = 24'b100110011001100110011001;
rgb[4874] = 24'b101010101010101010101010;
rgb[4875] = 24'b101110111011101110111011;
rgb[4876] = 24'b110011001100110011001100;
rgb[4877] = 24'b110111011101110111011101;
rgb[4878] = 24'b111011101110111011101110;
rgb[4879] = 24'b111111111111111111111111;
rgb[4880] = 24'b000000000000000000000000;
rgb[4881] = 24'b000100000001001000001111;
rgb[4882] = 24'b001000000010010000011111;
rgb[4883] = 24'b001100000011011000101111;
rgb[4884] = 24'b010000010100100000111111;
rgb[4885] = 24'b010100010101101001001111;
rgb[4886] = 24'b011000010110110001011111;
rgb[4887] = 24'b011100100111111001101111;
rgb[4888] = 24'b100000111000111110000000;
rgb[4889] = 24'b100101001001111110010010;
rgb[4890] = 24'b101001101010111110100100;
rgb[4891] = 24'b101110001011111110110110;
rgb[4892] = 24'b110010011100111111001000;
rgb[4893] = 24'b110110111101111111011010;
rgb[4894] = 24'b111011011110111111101100;
rgb[4895] = 24'b111111111111111111111111;
rgb[4896] = 24'b000000000000000000000000;
rgb[4897] = 24'b000011110001001100001110;
rgb[4898] = 24'b000111110010011000011101;
rgb[4899] = 24'b001011100011100100101100;
rgb[4900] = 24'b001111100100110100111010;
rgb[4901] = 24'b010011010110000001001001;
rgb[4902] = 24'b010111010111001101011000;
rgb[4903] = 24'b011011011000011001100111;
rgb[4904] = 24'b011111101001011101111000;
rgb[4905] = 24'b100100001010011010001011;
rgb[4906] = 24'b101000101011010110011110;
rgb[4907] = 24'b101101011100010010110001;
rgb[4908] = 24'b110001111101001011000101;
rgb[4909] = 24'b110110101110000111011000;
rgb[4910] = 24'b111011001111000011101011;
rgb[4911] = 24'b111111111111111111111111;
rgb[4912] = 24'b000000000000000000000000;
rgb[4913] = 24'b000011100001010000001101;
rgb[4914] = 24'b000111010010100000011011;
rgb[4915] = 24'b001011000011110100101000;
rgb[4916] = 24'b001110110101000100110110;
rgb[4917] = 24'b010010100110010101000100;
rgb[4918] = 24'b010110010111101001010001;
rgb[4919] = 24'b011010001000111001011111;
rgb[4920] = 24'b011110011001111101110000;
rgb[4921] = 24'b100011001010110110000100;
rgb[4922] = 24'b100111111011101110011000;
rgb[4923] = 24'b101100101100100010101101;
rgb[4924] = 24'b110001011101011011000001;
rgb[4925] = 24'b110110001110001111010110;
rgb[4926] = 24'b111010111111000111101010;
rgb[4927] = 24'b111111111111111111111111;
rgb[4928] = 24'b000000000000000000000000;
rgb[4929] = 24'b000011100001010100001100;
rgb[4930] = 24'b000111000010101100011000;
rgb[4931] = 24'b001010100100000000100101;
rgb[4932] = 24'b001110000101011000110001;
rgb[4933] = 24'b010001100110101100111110;
rgb[4934] = 24'b010101011000000101001010;
rgb[4935] = 24'b011000111001011001010111;
rgb[4936] = 24'b011101001010011101101000;
rgb[4937] = 24'b100010001011010001111101;
rgb[4938] = 24'b100110111100000010010011;
rgb[4939] = 24'b101011111100110110101000;
rgb[4940] = 24'b110000111101100110111110;
rgb[4941] = 24'b110101111110011011010011;
rgb[4942] = 24'b111010111111001011101001;
rgb[4943] = 24'b111111111111111111111111;
rgb[4944] = 24'b000000000000000000000000;
rgb[4945] = 24'b000011010001011000001011;
rgb[4946] = 24'b000110100010110100010110;
rgb[4947] = 24'b001010000100010000100010;
rgb[4948] = 24'b001101010101101000101101;
rgb[4949] = 24'b010000110111000100111000;
rgb[4950] = 24'b010100001000100001000100;
rgb[4951] = 24'b010111101001111001001111;
rgb[4952] = 24'b011011111010111101100000;
rgb[4953] = 24'b100000111011101101110110;
rgb[4954] = 24'b100110001100011010001101;
rgb[4955] = 24'b101011001101000110100100;
rgb[4956] = 24'b110000011101110110111011;
rgb[4957] = 24'b110101011110100011010001;
rgb[4958] = 24'b111010101111001111101000;
rgb[4959] = 24'b111111111111111111111111;
rgb[4960] = 24'b000000000000000000000000;
rgb[4961] = 24'b000011000001011100001010;
rgb[4962] = 24'b000110010010111100010100;
rgb[4963] = 24'b001001100100011100011110;
rgb[4964] = 24'b001100110101111100101000;
rgb[4965] = 24'b001111110111011000110011;
rgb[4966] = 24'b010011001000111000111101;
rgb[4967] = 24'b010110011010011001000111;
rgb[4968] = 24'b011010101011011101011000;
rgb[4969] = 24'b011111111100000101110000;
rgb[4970] = 24'b100101001100110010000111;
rgb[4971] = 24'b101010101101011010011111;
rgb[4972] = 24'b101111111110000010110111;
rgb[4973] = 24'b110101001110101011001111;
rgb[4974] = 24'b111010011111010011100111;
rgb[4975] = 24'b111111111111111011111111;
rgb[4976] = 24'b000000000000000000000000;
rgb[4977] = 24'b000011000001100000001001;
rgb[4978] = 24'b000110000011000100010010;
rgb[4979] = 24'b001001000100101000011011;
rgb[4980] = 24'b001100000110001100100100;
rgb[4981] = 24'b001111000111110000101101;
rgb[4982] = 24'b010010001001010100110110;
rgb[4983] = 24'b010101001010111000111111;
rgb[4984] = 24'b011001011011111101010000;
rgb[4985] = 24'b011110111100100001101001;
rgb[4986] = 24'b100100011101000110000010;
rgb[4987] = 24'b101001111101101010011011;
rgb[4988] = 24'b101111011110001110110100;
rgb[4989] = 24'b110100111110110011001101;
rgb[4990] = 24'b111010011111010111100110;
rgb[4991] = 24'b111111111111111111111111;
rgb[4992] = 24'b000000000000000000000000;
rgb[4993] = 24'b000010110001101000000111;
rgb[4994] = 24'b000101100011010000001111;
rgb[4995] = 24'b001000100100111000010111;
rgb[4996] = 24'b001011010110100000011111;
rgb[4997] = 24'b001110001000001000100111;
rgb[4998] = 24'b010001001001110000101111;
rgb[4999] = 24'b010011111011011000110111;
rgb[5000] = 24'b011000001100011101001000;
rgb[5001] = 24'b011101111100111101100010;
rgb[5002] = 24'b100011011101011101111100;
rgb[5003] = 24'b101001001101111110010110;
rgb[5004] = 24'b101110111110011110110000;
rgb[5005] = 24'b110100011110111111001010;
rgb[5006] = 24'b111010001111011111100100;
rgb[5007] = 24'b111111111111111011111111;
rgb[5008] = 24'b000000000000000000000000;
rgb[5009] = 24'b000010100001101100000110;
rgb[5010] = 24'b000101010011011000001101;
rgb[5011] = 24'b001000000101000100010100;
rgb[5012] = 24'b001010100110110000011011;
rgb[5013] = 24'b001101011000100000100001;
rgb[5014] = 24'b010000001010001100101000;
rgb[5015] = 24'b010010101011111000101111;
rgb[5016] = 24'b010110111100111101000000;
rgb[5017] = 24'b011100111101011001011011;
rgb[5018] = 24'b100010101101110101110110;
rgb[5019] = 24'b101000011110001110010010;
rgb[5020] = 24'b101110011110101010101101;
rgb[5021] = 24'b110100001111000111001000;
rgb[5022] = 24'b111001111111100011100011;
rgb[5023] = 24'b111111111111111111111111;
rgb[5024] = 24'b000000000000000000000000;
rgb[5025] = 24'b000010010001110000000101;
rgb[5026] = 24'b000100110011100000001011;
rgb[5027] = 24'b000111010101010100010001;
rgb[5028] = 24'b001001110111000100010110;
rgb[5029] = 24'b001100011000110100011100;
rgb[5030] = 24'b001110111010101000100010;
rgb[5031] = 24'b010001011100011000100111;
rgb[5032] = 24'b010101101101011100111000;
rgb[5033] = 24'b011011101101110101010100;
rgb[5034] = 24'b100001101110001001110001;
rgb[5035] = 24'b100111101110100010001101;
rgb[5036] = 24'b101101101110111010101010;
rgb[5037] = 24'b110011101111001111000110;
rgb[5038] = 24'b111001101111100111100010;
rgb[5039] = 24'b111111111111111011111111;
rgb[5040] = 24'b000000000000000000000000;
rgb[5041] = 24'b000010010001110100000100;
rgb[5042] = 24'b000100100011101000001001;
rgb[5043] = 24'b000110110101100000001101;
rgb[5044] = 24'b001001010111010100010010;
rgb[5045] = 24'b001011101001001100010110;
rgb[5046] = 24'b001101111011000000011011;
rgb[5047] = 24'b010000001100111000011111;
rgb[5048] = 24'b010100011101111100110000;
rgb[5049] = 24'b011010101110001101001110;
rgb[5050] = 24'b100000111110100001101011;
rgb[5051] = 24'b100111001110110010001001;
rgb[5052] = 24'b101101001111000110100110;
rgb[5053] = 24'b110011011111010111000100;
rgb[5054] = 24'b111001101111101011100001;
rgb[5055] = 24'b111111111111111111111111;
rgb[5056] = 24'b000000000000000000000000;
rgb[5057] = 24'b000010000001111000000011;
rgb[5058] = 24'b000100010011110100000110;
rgb[5059] = 24'b000110010101101100001010;
rgb[5060] = 24'b001000100111101000001101;
rgb[5061] = 24'b001010101001100100010000;
rgb[5062] = 24'b001100111011011100010100;
rgb[5063] = 24'b001111001101011000010111;
rgb[5064] = 24'b010011011110011100101000;
rgb[5065] = 24'b011001101110101001000111;
rgb[5066] = 24'b011111111110111001100101;
rgb[5067] = 24'b100110011111000110000100;
rgb[5068] = 24'b101100101111010010100011;
rgb[5069] = 24'b110011001111100011000001;
rgb[5070] = 24'b111001011111101111100000;
rgb[5071] = 24'b111111111111111111111111;
rgb[5072] = 24'b000000000000000000000000;
rgb[5073] = 24'b000001110001111100000010;
rgb[5074] = 24'b000011110011111100000100;
rgb[5075] = 24'b000101110101111100000110;
rgb[5076] = 24'b000111110111111000001001;
rgb[5077] = 24'b001001111001111000001011;
rgb[5078] = 24'b001011111011111000001101;
rgb[5079] = 24'b001101111101111000001111;
rgb[5080] = 24'b010010001110111100100000;
rgb[5081] = 24'b011000101111000101000000;
rgb[5082] = 24'b011111001111001101100000;
rgb[5083] = 24'b100101101111010110000000;
rgb[5084] = 24'b101100001111100010011111;
rgb[5085] = 24'b110010101111101010111111;
rgb[5086] = 24'b111001001111110011011111;
rgb[5087] = 24'b111111111111111111111111;
rgb[5088] = 24'b000000000000000000000000;
rgb[5089] = 24'b000001110010000000000001;
rgb[5090] = 24'b000011100100000100000010;
rgb[5091] = 24'b000101010110001000000011;
rgb[5092] = 24'b000111001000001100000100;
rgb[5093] = 24'b001000111010010000000101;
rgb[5094] = 24'b001010111100010100000110;
rgb[5095] = 24'b001100101110011000000111;
rgb[5096] = 24'b010000111111011100011000;
rgb[5097] = 24'b010111101111100000111001;
rgb[5098] = 24'b011110001111100101011010;
rgb[5099] = 24'b100100111111101001111011;
rgb[5100] = 24'b101011101111101110011100;
rgb[5101] = 24'b110010011111110010111101;
rgb[5102] = 24'b111001001111110111011110;
rgb[5103] = 24'b111111111111111111111111;
rgb[5104] = 24'b000000000000000000000000;
rgb[5105] = 24'b000001100010001000000000;
rgb[5106] = 24'b000011000100010000000000;
rgb[5107] = 24'b000100110110011000000000;
rgb[5108] = 24'b000110011000100000000000;
rgb[5109] = 24'b001000001010101000000000;
rgb[5110] = 24'b001001101100110000000000;
rgb[5111] = 24'b001011011110111000000000;
rgb[5112] = 24'b001111101111111000010001;
rgb[5113] = 24'b010110011111111100110010;
rgb[5114] = 24'b011101011111111001010101;
rgb[5115] = 24'b100100001111111101110110;
rgb[5116] = 24'b101011001111111110011001;
rgb[5117] = 24'b110001111111111110111011;
rgb[5118] = 24'b111000111111111111011101;
rgb[5119] = 24'b111111111111111111111111;
rgb[5120] = 24'b000000000000000000000000;
rgb[5121] = 24'b000100010001000100010001;
rgb[5122] = 24'b001000100010001000100010;
rgb[5123] = 24'b001100110011001100110011;
rgb[5124] = 24'b010001000100010001000100;
rgb[5125] = 24'b010101010101010101010101;
rgb[5126] = 24'b011001100110011001100110;
rgb[5127] = 24'b011101110111011101110111;
rgb[5128] = 24'b100010001000100010001000;
rgb[5129] = 24'b100110011001100110011001;
rgb[5130] = 24'b101010101010101010101010;
rgb[5131] = 24'b101110111011101110111011;
rgb[5132] = 24'b110011001100110011001100;
rgb[5133] = 24'b110111011101110111011101;
rgb[5134] = 24'b111011101110111011101110;
rgb[5135] = 24'b111111111111111111111111;
rgb[5136] = 24'b000000000000000000000000;
rgb[5137] = 24'b000100000001001000001111;
rgb[5138] = 24'b001000000010010000011111;
rgb[5139] = 24'b001100000011011000101111;
rgb[5140] = 24'b010000000100100000111111;
rgb[5141] = 24'b010100000101101001001111;
rgb[5142] = 24'b011000000110110001011111;
rgb[5143] = 24'b011100000111111001101111;
rgb[5144] = 24'b100000011000111110000000;
rgb[5145] = 24'b100100111001111110010010;
rgb[5146] = 24'b101001011010111110100100;
rgb[5147] = 24'b101101111011111110110110;
rgb[5148] = 24'b110010011100111111001000;
rgb[5149] = 24'b110110111101111111011010;
rgb[5150] = 24'b111011011110111111101100;
rgb[5151] = 24'b111111111111111111111111;
rgb[5152] = 24'b000000000000000000000000;
rgb[5153] = 24'b000011110001001100001110;
rgb[5154] = 24'b000111100010011000011101;
rgb[5155] = 24'b001011010011100100101100;
rgb[5156] = 24'b001111000100110100111010;
rgb[5157] = 24'b010010110110000001001001;
rgb[5158] = 24'b010110100111001101011000;
rgb[5159] = 24'b011010101000011001100111;
rgb[5160] = 24'b011110111001011101111000;
rgb[5161] = 24'b100011011010011010001011;
rgb[5162] = 24'b101000001011010110011110;
rgb[5163] = 24'b101100111100010010110001;
rgb[5164] = 24'b110001101101001011000101;
rgb[5165] = 24'b110110011110000111011000;
rgb[5166] = 24'b111011001111000011101011;
rgb[5167] = 24'b111111111111111111111111;
rgb[5168] = 24'b000000000000000000000000;
rgb[5169] = 24'b000011100001010000001101;
rgb[5170] = 24'b000111000010100000011011;
rgb[5171] = 24'b001010100011110100101000;
rgb[5172] = 24'b001110000101000100110110;
rgb[5173] = 24'b010001110110010101000100;
rgb[5174] = 24'b010101010111101001010001;
rgb[5175] = 24'b011000111000111001011111;
rgb[5176] = 24'b011101001001111101110000;
rgb[5177] = 24'b100010001010110110000100;
rgb[5178] = 24'b100111001011101110011000;
rgb[5179] = 24'b101011111100100010101101;
rgb[5180] = 24'b110000111101011011000001;
rgb[5181] = 24'b110101111110001111010110;
rgb[5182] = 24'b111010111111000111101010;
rgb[5183] = 24'b111111111111111111111111;
rgb[5184] = 24'b000000000000000000000000;
rgb[5185] = 24'b000011010001010100001100;
rgb[5186] = 24'b000110100010101100011000;
rgb[5187] = 24'b001001110100000000100101;
rgb[5188] = 24'b001101010101011000110001;
rgb[5189] = 24'b010000100110101100111110;
rgb[5190] = 24'b010011111000000101001010;
rgb[5191] = 24'b010111011001011001010111;
rgb[5192] = 24'b011011101010011101101000;
rgb[5193] = 24'b100000101011010001111101;
rgb[5194] = 24'b100101111100000010010011;
rgb[5195] = 24'b101011001100110110101000;
rgb[5196] = 24'b110000001101100110111110;
rgb[5197] = 24'b110101011110011011010011;
rgb[5198] = 24'b111010101111001011101001;
rgb[5199] = 24'b111111111111111111111111;
rgb[5200] = 24'b000000000000000000000000;
rgb[5201] = 24'b000011000001011000001011;
rgb[5202] = 24'b000110000010110100010110;
rgb[5203] = 24'b001001010100010000100010;
rgb[5204] = 24'b001100010101101000101101;
rgb[5205] = 24'b001111100111000100111000;
rgb[5206] = 24'b010010101000100001000100;
rgb[5207] = 24'b010101101001111001001111;
rgb[5208] = 24'b011001111010111101100000;
rgb[5209] = 24'b011111011011101101110110;
rgb[5210] = 24'b100100111100011010001101;
rgb[5211] = 24'b101010001101000110100100;
rgb[5212] = 24'b101111101101110110111011;
rgb[5213] = 24'b110100111110100011010001;
rgb[5214] = 24'b111010011111001111101000;
rgb[5215] = 24'b111111111111111111111111;
rgb[5216] = 24'b000000000000000000000000;
rgb[5217] = 24'b000010110001011100001010;
rgb[5218] = 24'b000101100010111100010100;
rgb[5219] = 24'b001000100100011100011110;
rgb[5220] = 24'b001011010101111100101000;
rgb[5221] = 24'b001110010111011000110011;
rgb[5222] = 24'b010001001000111000111101;
rgb[5223] = 24'b010100001010011001000111;
rgb[5224] = 24'b011000011011011101011000;
rgb[5225] = 24'b011101111100000101110000;
rgb[5226] = 24'b100011101100110010000111;
rgb[5227] = 24'b101001001101011010011111;
rgb[5228] = 24'b101110111110000010110111;
rgb[5229] = 24'b110100011110101011001111;
rgb[5230] = 24'b111010001111010011100111;
rgb[5231] = 24'b111111111111111011111111;
rgb[5232] = 24'b000000000000000000000000;
rgb[5233] = 24'b000010100001100000001001;
rgb[5234] = 24'b000101010011000100010010;
rgb[5235] = 24'b000111110100101000011011;
rgb[5236] = 24'b001010100110001100100100;
rgb[5237] = 24'b001101000111110000101101;
rgb[5238] = 24'b001111111001010100110110;
rgb[5239] = 24'b010010101010111000111111;
rgb[5240] = 24'b010110111011111101010000;
rgb[5241] = 24'b011100101100100001101001;
rgb[5242] = 24'b100010011101000110000010;
rgb[5243] = 24'b101000011101101010011011;
rgb[5244] = 24'b101110001110001110110100;
rgb[5245] = 24'b110100001110110011001101;
rgb[5246] = 24'b111001111111010111100110;
rgb[5247] = 24'b111111111111111111111111;
rgb[5248] = 24'b000000000000000000000000;
rgb[5249] = 24'b000010010001101000000111;
rgb[5250] = 24'b000100110011010000001111;
rgb[5251] = 24'b000111000100111000010111;
rgb[5252] = 24'b001001100110100000011111;
rgb[5253] = 24'b001100001000001000100111;
rgb[5254] = 24'b001110011001110000101111;
rgb[5255] = 24'b010000111011011000110111;
rgb[5256] = 24'b010101001100011101001000;
rgb[5257] = 24'b011011001100111101100010;
rgb[5258] = 24'b100001011101011101111100;
rgb[5259] = 24'b100111011101111110010110;
rgb[5260] = 24'b101101011110011110110000;
rgb[5261] = 24'b110011101110111111001010;
rgb[5262] = 24'b111001101111011111100100;
rgb[5263] = 24'b111111111111111011111111;
rgb[5264] = 24'b000000000000000000000000;
rgb[5265] = 24'b000010000001101100000110;
rgb[5266] = 24'b000100010011011000001101;
rgb[5267] = 24'b000110100101000100010100;
rgb[5268] = 24'b001000100110110000011011;
rgb[5269] = 24'b001010111000100000100001;
rgb[5270] = 24'b001101001010001100101000;
rgb[5271] = 24'b001111011011111000101111;
rgb[5272] = 24'b010011101100111101000000;
rgb[5273] = 24'b011001111101011001011011;
rgb[5274] = 24'b100000001101110101110110;
rgb[5275] = 24'b100110011110001110010010;
rgb[5276] = 24'b101100111110101010101101;
rgb[5277] = 24'b110011001111000111001000;
rgb[5278] = 24'b111001011111100011100011;
rgb[5279] = 24'b111111111111111111111111;
rgb[5280] = 24'b000000000000000000000000;
rgb[5281] = 24'b000001110001110000000101;
rgb[5282] = 24'b000011110011100000001011;
rgb[5283] = 24'b000101110101010100010001;
rgb[5284] = 24'b000111110111000100010110;
rgb[5285] = 24'b001001111000110100011100;
rgb[5286] = 24'b001011101010101000100010;
rgb[5287] = 24'b001101101100011000100111;
rgb[5288] = 24'b010001111101011100111000;
rgb[5289] = 24'b011000011101110101010100;
rgb[5290] = 24'b011111001110001001110001;
rgb[5291] = 24'b100101101110100010001101;
rgb[5292] = 24'b101100001110111010101010;
rgb[5293] = 24'b110010101111001111000110;
rgb[5294] = 24'b111001001111100111100010;
rgb[5295] = 24'b111111111111111011111111;
rgb[5296] = 24'b000000000000000000000000;
rgb[5297] = 24'b000001100001110100000100;
rgb[5298] = 24'b000011010011101000001001;
rgb[5299] = 24'b000101000101100000001101;
rgb[5300] = 24'b000110110111010100010010;
rgb[5301] = 24'b001000101001001100010110;
rgb[5302] = 24'b001010011011000000011011;
rgb[5303] = 24'b001100001100111000011111;
rgb[5304] = 24'b010000011101111100110000;
rgb[5305] = 24'b010111001110001101001110;
rgb[5306] = 24'b011101111110100001101011;
rgb[5307] = 24'b100100101110110010001001;
rgb[5308] = 24'b101011011111000110100110;
rgb[5309] = 24'b110010001111010111000100;
rgb[5310] = 24'b111000111111101011100001;
rgb[5311] = 24'b111111111111111111111111;
rgb[5312] = 24'b000000000000000000000000;
rgb[5313] = 24'b000001010001111000000011;
rgb[5314] = 24'b000010110011110100000110;
rgb[5315] = 24'b000100010101101100001010;
rgb[5316] = 24'b000101110111101000001101;
rgb[5317] = 24'b000111011001100100010000;
rgb[5318] = 24'b001000111011011100010100;
rgb[5319] = 24'b001010011101011000010111;
rgb[5320] = 24'b001110101110011100101000;
rgb[5321] = 24'b010101101110101001000111;
rgb[5322] = 24'b011100101110111001100101;
rgb[5323] = 24'b100011101111000110000100;
rgb[5324] = 24'b101010101111010010100011;
rgb[5325] = 24'b110001101111100011000001;
rgb[5326] = 24'b111000101111101111100000;
rgb[5327] = 24'b111111111111111111111111;
rgb[5328] = 24'b000000000000000000000000;
rgb[5329] = 24'b000001010001111100000010;
rgb[5330] = 24'b000010100011111100000100;
rgb[5331] = 24'b000011110101111100000110;
rgb[5332] = 24'b000101000111111000001001;
rgb[5333] = 24'b000110011001111000001011;
rgb[5334] = 24'b000111101011111000001101;
rgb[5335] = 24'b001000111101111000001111;
rgb[5336] = 24'b001101001110111100100000;
rgb[5337] = 24'b010100011111000101000000;
rgb[5338] = 24'b011011101111001101100000;
rgb[5339] = 24'b100010111111010110000000;
rgb[5340] = 24'b101010001111100010011111;
rgb[5341] = 24'b110001011111101010111111;
rgb[5342] = 24'b111000101111110011011111;
rgb[5343] = 24'b111111111111111111111111;
rgb[5344] = 24'b000000000000000000000000;
rgb[5345] = 24'b000001000010000000000001;
rgb[5346] = 24'b000010000100000100000010;
rgb[5347] = 24'b000011000110001000000011;
rgb[5348] = 24'b000100001000001100000100;
rgb[5349] = 24'b000101001010010000000101;
rgb[5350] = 24'b000110001100010100000110;
rgb[5351] = 24'b000111011110011000000111;
rgb[5352] = 24'b001011101111011100011000;
rgb[5353] = 24'b010010111111100000111001;
rgb[5354] = 24'b011010011111100101011010;
rgb[5355] = 24'b100001111111101001111011;
rgb[5356] = 24'b101001011111101110011100;
rgb[5357] = 24'b110000111111110010111101;
rgb[5358] = 24'b111000011111110111011110;
rgb[5359] = 24'b111111111111111111111111;
rgb[5360] = 24'b000000000000000000000000;
rgb[5361] = 24'b000000110010001000000000;
rgb[5362] = 24'b000001100100010000000000;
rgb[5363] = 24'b000010010110011000000000;
rgb[5364] = 24'b000011001000100000000000;
rgb[5365] = 24'b000100001010101000000000;
rgb[5366] = 24'b000100111100110000000000;
rgb[5367] = 24'b000101101110111000000000;
rgb[5368] = 24'b001001111111111000010001;
rgb[5369] = 24'b010001101111111100110010;
rgb[5370] = 24'b011001011111111001010101;
rgb[5371] = 24'b100000111111111101110110;
rgb[5372] = 24'b101000101111111110011001;
rgb[5373] = 24'b110000011111111110111011;
rgb[5374] = 24'b111000001111111111011101;
rgb[5375] = 24'b111111111111111111111111;
rgb[5376] = 24'b000000000000000000000000;
rgb[5377] = 24'b000100010001000100010001;
rgb[5378] = 24'b001000100010001000100010;
rgb[5379] = 24'b001100110011001100110011;
rgb[5380] = 24'b010001000100010001000100;
rgb[5381] = 24'b010101010101010101010101;
rgb[5382] = 24'b011001100110011001100110;
rgb[5383] = 24'b011101110111011101110111;
rgb[5384] = 24'b100010001000100010001000;
rgb[5385] = 24'b100110011001100110011001;
rgb[5386] = 24'b101010101010101010101010;
rgb[5387] = 24'b101110111011101110111011;
rgb[5388] = 24'b110011001100110011001100;
rgb[5389] = 24'b110111011101110111011101;
rgb[5390] = 24'b111011101110111011101110;
rgb[5391] = 24'b111111111111111111111111;
rgb[5392] = 24'b000000000000000000000000;
rgb[5393] = 24'b000011110001001000001111;
rgb[5394] = 24'b000111110010010000011111;
rgb[5395] = 24'b001011110011011000101111;
rgb[5396] = 24'b001111110100100000111111;
rgb[5397] = 24'b010011110101101001001111;
rgb[5398] = 24'b010111110110110001011111;
rgb[5399] = 24'b011011110111111001101111;
rgb[5400] = 24'b100000001000111110000000;
rgb[5401] = 24'b100100101001111110010010;
rgb[5402] = 24'b101001001010111110100100;
rgb[5403] = 24'b101101101011111110110110;
rgb[5404] = 24'b110010001100111111001000;
rgb[5405] = 24'b110110101101111111011010;
rgb[5406] = 24'b111011001110111111101100;
rgb[5407] = 24'b111111111111111111111111;
rgb[5408] = 24'b000000000000000000000000;
rgb[5409] = 24'b000011100001001100001110;
rgb[5410] = 24'b000111010010011000011101;
rgb[5411] = 24'b001011000011100100101100;
rgb[5412] = 24'b001110100100110100111010;
rgb[5413] = 24'b010010010110000001001001;
rgb[5414] = 24'b010110000111001101011000;
rgb[5415] = 24'b011001111000011001100111;
rgb[5416] = 24'b011110001001011101111000;
rgb[5417] = 24'b100010111010011010001011;
rgb[5418] = 24'b100111101011010110011110;
rgb[5419] = 24'b101100011100010010110001;
rgb[5420] = 24'b110001011101001011000101;
rgb[5421] = 24'b110110001110000111011000;
rgb[5422] = 24'b111010111111000011101011;
rgb[5423] = 24'b111111111111111111111111;
rgb[5424] = 24'b000000000000000000000000;
rgb[5425] = 24'b000011010001010000001101;
rgb[5426] = 24'b000110110010100000011011;
rgb[5427] = 24'b001010000011110100101000;
rgb[5428] = 24'b001101100101000100110110;
rgb[5429] = 24'b010001000110010101000100;
rgb[5430] = 24'b010100010111101001010001;
rgb[5431] = 24'b010111111000111001011111;
rgb[5432] = 24'b011100001001111101110000;
rgb[5433] = 24'b100001001010110110000100;
rgb[5434] = 24'b100110001011101110011000;
rgb[5435] = 24'b101011011100100010101101;
rgb[5436] = 24'b110000011101011011000001;
rgb[5437] = 24'b110101101110001111010110;
rgb[5438] = 24'b111010101111000111101010;
rgb[5439] = 24'b111111111111111111111111;
rgb[5440] = 24'b000000000000000000000000;
rgb[5441] = 24'b000011000001010100001100;
rgb[5442] = 24'b000110000010101100011000;
rgb[5443] = 24'b001001010100000000100101;
rgb[5444] = 24'b001100010101011000110001;
rgb[5445] = 24'b001111100110101100111110;
rgb[5446] = 24'b010010101000000101001010;
rgb[5447] = 24'b010101111001011001010111;
rgb[5448] = 24'b011010001010011101101000;
rgb[5449] = 24'b011111011011010001111101;
rgb[5450] = 24'b100100111100000010010011;
rgb[5451] = 24'b101010001100110110101000;
rgb[5452] = 24'b101111101101100110111110;
rgb[5453] = 24'b110100111110011011010011;
rgb[5454] = 24'b111010011111001011101001;
rgb[5455] = 24'b111111111111111111111111;
rgb[5456] = 24'b000000000000000000000000;
rgb[5457] = 24'b000010110001011000001011;
rgb[5458] = 24'b000101100010110100010110;
rgb[5459] = 24'b001000100100010000100010;
rgb[5460] = 24'b001011010101101000101101;
rgb[5461] = 24'b001110000111000100111000;
rgb[5462] = 24'b010001001000100001000100;
rgb[5463] = 24'b010011111001111001001111;
rgb[5464] = 24'b011000001010111101100000;
rgb[5465] = 24'b011101101011101101110110;
rgb[5466] = 24'b100011011100011010001101;
rgb[5467] = 24'b101001001101000110100100;
rgb[5468] = 24'b101110111101110110111011;
rgb[5469] = 24'b110100011110100011010001;
rgb[5470] = 24'b111010001111001111101000;
rgb[5471] = 24'b111111111111111111111111;
rgb[5472] = 24'b000000000000000000000000;
rgb[5473] = 24'b000010100001011100001010;
rgb[5474] = 24'b000101000010111100010100;
rgb[5475] = 24'b000111100100011100011110;
rgb[5476] = 24'b001010000101111100101000;
rgb[5477] = 24'b001100110111011000110011;
rgb[5478] = 24'b001111011000111000111101;
rgb[5479] = 24'b010001111010011001000111;
rgb[5480] = 24'b010110001011011101011000;
rgb[5481] = 24'b011100001100000101110000;
rgb[5482] = 24'b100001111100110010000111;
rgb[5483] = 24'b100111111101011010011111;
rgb[5484] = 24'b101101111110000010110111;
rgb[5485] = 24'b110011111110101011001111;
rgb[5486] = 24'b111001111111010011100111;
rgb[5487] = 24'b111111111111111011111111;
rgb[5488] = 24'b000000000000000000000000;
rgb[5489] = 24'b000010010001100000001001;
rgb[5490] = 24'b000100100011000100010010;
rgb[5491] = 24'b000110110100101000011011;
rgb[5492] = 24'b001001000110001100100100;
rgb[5493] = 24'b001011010111110000101101;
rgb[5494] = 24'b001101101001010100110110;
rgb[5495] = 24'b001111111010111000111111;
rgb[5496] = 24'b010100001011111101010000;
rgb[5497] = 24'b011010011100100001101001;
rgb[5498] = 24'b100000101101000110000010;
rgb[5499] = 24'b100110111101101010011011;
rgb[5500] = 24'b101101001110001110110100;
rgb[5501] = 24'b110011011110110011001101;
rgb[5502] = 24'b111001101111010111100110;
rgb[5503] = 24'b111111111111111111111111;
rgb[5504] = 24'b000000000000000000000000;
rgb[5505] = 24'b000001110001101000000111;
rgb[5506] = 24'b000011110011010000001111;
rgb[5507] = 24'b000101110100111000010111;
rgb[5508] = 24'b000111110110100000011111;
rgb[5509] = 24'b001001111000001000100111;
rgb[5510] = 24'b001011111001110000101111;
rgb[5511] = 24'b001101111011011000110111;
rgb[5512] = 24'b010010001100011101001000;
rgb[5513] = 24'b011000101100111101100010;
rgb[5514] = 24'b011111001101011101111100;
rgb[5515] = 24'b100101101101111110010110;
rgb[5516] = 24'b101100001110011110110000;
rgb[5517] = 24'b110010101110111111001010;
rgb[5518] = 24'b111001001111011111100100;
rgb[5519] = 24'b111111111111111011111111;
rgb[5520] = 24'b000000000000000000000000;
rgb[5521] = 24'b000001100001101100000110;
rgb[5522] = 24'b000011010011011000001101;
rgb[5523] = 24'b000101000101000100010100;
rgb[5524] = 24'b000110110110110000011011;
rgb[5525] = 24'b001000011000100000100001;
rgb[5526] = 24'b001010001010001100101000;
rgb[5527] = 24'b001011111011111000101111;
rgb[5528] = 24'b010000001100111101000000;
rgb[5529] = 24'b010110111101011001011011;
rgb[5530] = 24'b011101101101110101110110;
rgb[5531] = 24'b100100101110001110010010;
rgb[5532] = 24'b101011011110101010101101;
rgb[5533] = 24'b110010001111000111001000;
rgb[5534] = 24'b111000111111100011100011;
rgb[5535] = 24'b111111111111111111111111;
rgb[5536] = 24'b000000000000000000000000;
rgb[5537] = 24'b000001010001110000000101;
rgb[5538] = 24'b000010110011100000001011;
rgb[5539] = 24'b000100010101010100010001;
rgb[5540] = 24'b000101100111000100010110;
rgb[5541] = 24'b000111001000110100011100;
rgb[5542] = 24'b001000101010101000100010;
rgb[5543] = 24'b001001111100011000100111;
rgb[5544] = 24'b001110001101011100111000;
rgb[5545] = 24'b010101001101110101010100;
rgb[5546] = 24'b011100011110001001110001;
rgb[5547] = 24'b100011011110100010001101;
rgb[5548] = 24'b101010101110111010101010;
rgb[5549] = 24'b110001101111001111000110;
rgb[5550] = 24'b111000101111100111100010;
rgb[5551] = 24'b111111111111111011111111;
rgb[5552] = 24'b000000000000000000000000;
rgb[5553] = 24'b000001000001110100000100;
rgb[5554] = 24'b000010010011101000001001;
rgb[5555] = 24'b000011010101100000001101;
rgb[5556] = 24'b000100100111010100010010;
rgb[5557] = 24'b000101101001001100010110;
rgb[5558] = 24'b000110111011000000011011;
rgb[5559] = 24'b000111111100111000011111;
rgb[5560] = 24'b001100001101111100110000;
rgb[5561] = 24'b010011101110001101001110;
rgb[5562] = 24'b011010111110100001101011;
rgb[5563] = 24'b100010011110110010001001;
rgb[5564] = 24'b101001101111000110100110;
rgb[5565] = 24'b110001001111010111000100;
rgb[5566] = 24'b111000011111101011100001;
rgb[5567] = 24'b111111111111111111111111;
rgb[5568] = 24'b000000000000000000000000;
rgb[5569] = 24'b000000110001111000000011;
rgb[5570] = 24'b000001100011110100000110;
rgb[5571] = 24'b000010100101101100001010;
rgb[5572] = 24'b000011010111101000001101;
rgb[5573] = 24'b000100001001100100010000;
rgb[5574] = 24'b000101001011011100010100;
rgb[5575] = 24'b000101111101011000010111;
rgb[5576] = 24'b001010001110011100101000;
rgb[5577] = 24'b010001111110101001000111;
rgb[5578] = 24'b011001011110111001100101;
rgb[5579] = 24'b100001001111000110000100;
rgb[5580] = 24'b101000111111010010100011;
rgb[5581] = 24'b110000011111100011000001;
rgb[5582] = 24'b111000001111101111100000;
rgb[5583] = 24'b111111111111111111111111;
rgb[5584] = 24'b000000000000000000000000;
rgb[5585] = 24'b000000100001111100000010;
rgb[5586] = 24'b000001000011111100000100;
rgb[5587] = 24'b000001100101111100000110;
rgb[5588] = 24'b000010010111111000001001;
rgb[5589] = 24'b000010111001111000001011;
rgb[5590] = 24'b000011011011111000001101;
rgb[5591] = 24'b000011111101111000001111;
rgb[5592] = 24'b001000001110111100100000;
rgb[5593] = 24'b010000001111000101000000;
rgb[5594] = 24'b011000001111001101100000;
rgb[5595] = 24'b100000001111010110000000;
rgb[5596] = 24'b100111111111100010011111;
rgb[5597] = 24'b101111111111101010111111;
rgb[5598] = 24'b110111111111110011011111;
rgb[5599] = 24'b111111111111111111111111;
rgb[5600] = 24'b000000000000000000000000;
rgb[5601] = 24'b000000010010000000000001;
rgb[5602] = 24'b000000100100000100000010;
rgb[5603] = 24'b000000110110001000000011;
rgb[5604] = 24'b000001001000001100000100;
rgb[5605] = 24'b000001011010010000000101;
rgb[5606] = 24'b000001101100010100000110;
rgb[5607] = 24'b000001111110011000000111;
rgb[5608] = 24'b000110001111011100011000;
rgb[5609] = 24'b001110011111100000111001;
rgb[5610] = 24'b010110101111100101011010;
rgb[5611] = 24'b011110111111101001111011;
rgb[5612] = 24'b100111001111101110011100;
rgb[5613] = 24'b101111011111110010111101;
rgb[5614] = 24'b110111101111110111011110;
rgb[5615] = 24'b111111111111111111111111;
rgb[5616] = 24'b000000000000000000000000;
rgb[5617] = 24'b000000000010001000000000;
rgb[5618] = 24'b000000000100010000000000;
rgb[5619] = 24'b000000000110011000000000;
rgb[5620] = 24'b000000001000100000000000;
rgb[5621] = 24'b000000001010101000000000;
rgb[5622] = 24'b000000001100110000000000;
rgb[5623] = 24'b000000001110111000000000;
rgb[5624] = 24'b000100011111111000010001;
rgb[5625] = 24'b001100101111111100110010;
rgb[5626] = 24'b010101011111111001010101;
rgb[5627] = 24'b011101101111111101110110;
rgb[5628] = 24'b100110011111111110011001;
rgb[5629] = 24'b101110111111111110111011;
rgb[5630] = 24'b110111011111111111011101;
rgb[5631] = 24'b111111111111111111111111;
rgb[5632] = 24'b000000000000000000000000;
rgb[5633] = 24'b000100010001000100010001;
rgb[5634] = 24'b001000100010001000100010;
rgb[5635] = 24'b001100110011001100110011;
rgb[5636] = 24'b010001000100010001000100;
rgb[5637] = 24'b010101010101010101010101;
rgb[5638] = 24'b011001100110011001100110;
rgb[5639] = 24'b011101110111011101110111;
rgb[5640] = 24'b100010001000100010001000;
rgb[5641] = 24'b100110011001100110011001;
rgb[5642] = 24'b101010101010101010101010;
rgb[5643] = 24'b101110111011101110111011;
rgb[5644] = 24'b110011001100110011001100;
rgb[5645] = 24'b110111011101110111011101;
rgb[5646] = 24'b111011101110111011101110;
rgb[5647] = 24'b111111111111111111111111;
rgb[5648] = 24'b000000000000000000000000;
rgb[5649] = 24'b000011110001001000010000;
rgb[5650] = 24'b000111110010010000100000;
rgb[5651] = 24'b001011110011011000110000;
rgb[5652] = 24'b001111110100100001000000;
rgb[5653] = 24'b010011110101101001010000;
rgb[5654] = 24'b010111110110110001100000;
rgb[5655] = 24'b011011110111111001110000;
rgb[5656] = 24'b100000001000111110000001;
rgb[5657] = 24'b100100101001111110010011;
rgb[5658] = 24'b101001001010111110100101;
rgb[5659] = 24'b101101101011111110110111;
rgb[5660] = 24'b110010001100111111001001;
rgb[5661] = 24'b110110101101111111011011;
rgb[5662] = 24'b111011001110111111101101;
rgb[5663] = 24'b111111111111111111111111;
rgb[5664] = 24'b000000000000000000000000;
rgb[5665] = 24'b000011100001001100001111;
rgb[5666] = 24'b000111010010011000011110;
rgb[5667] = 24'b001011000011100100101101;
rgb[5668] = 24'b001110100100110100111100;
rgb[5669] = 24'b010010010110000001001011;
rgb[5670] = 24'b010110000111001101011010;
rgb[5671] = 24'b011001111000011001101010;
rgb[5672] = 24'b011110001001011101111011;
rgb[5673] = 24'b100010111010011010001101;
rgb[5674] = 24'b100111101011010110100000;
rgb[5675] = 24'b101100011100010010110011;
rgb[5676] = 24'b110001011101001011000110;
rgb[5677] = 24'b110110001110000111011001;
rgb[5678] = 24'b111010111111000011101100;
rgb[5679] = 24'b111111111111111111111111;
rgb[5680] = 24'b000000000000000000000000;
rgb[5681] = 24'b000011010001010000001110;
rgb[5682] = 24'b000110110010100000011100;
rgb[5683] = 24'b001010000011110100101010;
rgb[5684] = 24'b001101100101000100111000;
rgb[5685] = 24'b010001000110010101000111;
rgb[5686] = 24'b010100010111101001010101;
rgb[5687] = 24'b010111111000111001100011;
rgb[5688] = 24'b011100001001111101110100;
rgb[5689] = 24'b100001001010110110001000;
rgb[5690] = 24'b100110001011101110011100;
rgb[5691] = 24'b101011011100100010101111;
rgb[5692] = 24'b110000011101011011000011;
rgb[5693] = 24'b110101101110001111010111;
rgb[5694] = 24'b111010101111000111101011;
rgb[5695] = 24'b111111111111111111111111;
rgb[5696] = 24'b000000000000000000000000;
rgb[5697] = 24'b000011000001010100001101;
rgb[5698] = 24'b000110000010101100011010;
rgb[5699] = 24'b001001010100000000100111;
rgb[5700] = 24'b001100010101011000110101;
rgb[5701] = 24'b001111100110101101000010;
rgb[5702] = 24'b010010101000000101001111;
rgb[5703] = 24'b010101111001011001011101;
rgb[5704] = 24'b011010001010011101101110;
rgb[5705] = 24'b011111011011010010000010;
rgb[5706] = 24'b100100111100000010010111;
rgb[5707] = 24'b101010001100110110101100;
rgb[5708] = 24'b101111101101100111000000;
rgb[5709] = 24'b110100111110011011010101;
rgb[5710] = 24'b111010011111001011101010;
rgb[5711] = 24'b111111111111111111111111;
rgb[5712] = 24'b000000000000000000000000;
rgb[5713] = 24'b000010110001011000001100;
rgb[5714] = 24'b000101100010110100011000;
rgb[5715] = 24'b001000100100010000100101;
rgb[5716] = 24'b001011010101101000110001;
rgb[5717] = 24'b001110000111000100111110;
rgb[5718] = 24'b010001001000100001001010;
rgb[5719] = 24'b010011111001111001010110;
rgb[5720] = 24'b011000001010111101100111;
rgb[5721] = 24'b011101101011101101111101;
rgb[5722] = 24'b100011011100011010010011;
rgb[5723] = 24'b101001001101000110101000;
rgb[5724] = 24'b101110111101110110111110;
rgb[5725] = 24'b110100011110100011010011;
rgb[5726] = 24'b111010001111001111101001;
rgb[5727] = 24'b111111111111111111111111;
rgb[5728] = 24'b000000000000000000000000;
rgb[5729] = 24'b000010100001011100001011;
rgb[5730] = 24'b000101000010111100010110;
rgb[5731] = 24'b000111100100011100100010;
rgb[5732] = 24'b001010000101111100101101;
rgb[5733] = 24'b001100110111011000111001;
rgb[5734] = 24'b001111011000111001000100;
rgb[5735] = 24'b010001111010011001010000;
rgb[5736] = 24'b010110001011011101100001;
rgb[5737] = 24'b011100001100000101110111;
rgb[5738] = 24'b100001111100110010001110;
rgb[5739] = 24'b100111111101011010100100;
rgb[5740] = 24'b101101111110000010111011;
rgb[5741] = 24'b110011111110101011010001;
rgb[5742] = 24'b111001111111010011101000;
rgb[5743] = 24'b111111111111111011111111;
rgb[5744] = 24'b000000000000000000000000;
rgb[5745] = 24'b000010010001100000001010;
rgb[5746] = 24'b000100100011000100010101;
rgb[5747] = 24'b000110110100101000011111;
rgb[5748] = 24'b001001000110001100101010;
rgb[5749] = 24'b001011010111110000110100;
rgb[5750] = 24'b001101101001010100111111;
rgb[5751] = 24'b001111111010111001001010;
rgb[5752] = 24'b010100001011111101011011;
rgb[5753] = 24'b011010011100100001110010;
rgb[5754] = 24'b100000101101000110001001;
rgb[5755] = 24'b100110111101101010100001;
rgb[5756] = 24'b101101001110001110111000;
rgb[5757] = 24'b110011011110110011010000;
rgb[5758] = 24'b111001101111010111100111;
rgb[5759] = 24'b111111111111111111111111;
rgb[5760] = 24'b000000000000000000000000;
rgb[5761] = 24'b000001110001101000001001;
rgb[5762] = 24'b000011110011010000010011;
rgb[5763] = 24'b000101110100111000011100;
rgb[5764] = 24'b000111110110100000100110;
rgb[5765] = 24'b001001111000001000110000;
rgb[5766] = 24'b001011111001110000111001;
rgb[5767] = 24'b001101111011011001000011;
rgb[5768] = 24'b010010001100011101010100;
rgb[5769] = 24'b011000101100111101101100;
rgb[5770] = 24'b011111001101011110000101;
rgb[5771] = 24'b100101101101111110011101;
rgb[5772] = 24'b101100001110011110110101;
rgb[5773] = 24'b110010101110111111001110;
rgb[5774] = 24'b111001001111011111100110;
rgb[5775] = 24'b111111111111111011111111;
rgb[5776] = 24'b000000000000000000000000;
rgb[5777] = 24'b000001100001101100001000;
rgb[5778] = 24'b000011010011011000010001;
rgb[5779] = 24'b000101000101000100011010;
rgb[5780] = 24'b000110110110110000100010;
rgb[5781] = 24'b001000011000100000101011;
rgb[5782] = 24'b001010001010001100110100;
rgb[5783] = 24'b001011111011111000111101;
rgb[5784] = 24'b010000001100111101001110;
rgb[5785] = 24'b010110111101011001100111;
rgb[5786] = 24'b011101101101110110000000;
rgb[5787] = 24'b100100101110001110011001;
rgb[5788] = 24'b101011011110101010110011;
rgb[5789] = 24'b110010001111000111001100;
rgb[5790] = 24'b111000111111100011100101;
rgb[5791] = 24'b111111111111111111111111;
rgb[5792] = 24'b000000000000000000000000;
rgb[5793] = 24'b000001010001110000000111;
rgb[5794] = 24'b000010110011100000001111;
rgb[5795] = 24'b000100010101010100010111;
rgb[5796] = 24'b000101100111000100011111;
rgb[5797] = 24'b000111001000110100100111;
rgb[5798] = 24'b001000101010101000101110;
rgb[5799] = 24'b001001111100011000110110;
rgb[5800] = 24'b001110001101011101000111;
rgb[5801] = 24'b010101001101110101100001;
rgb[5802] = 24'b011100011110001001111100;
rgb[5803] = 24'b100011011110100010010110;
rgb[5804] = 24'b101010101110111010110000;
rgb[5805] = 24'b110001101111001111001010;
rgb[5806] = 24'b111000101111100111100100;
rgb[5807] = 24'b111111111111111011111111;
rgb[5808] = 24'b000000000000000000000000;
rgb[5809] = 24'b000001000001110100000110;
rgb[5810] = 24'b000010010011101000001101;
rgb[5811] = 24'b000011010101100000010100;
rgb[5812] = 24'b000100100111010100011011;
rgb[5813] = 24'b000101101001001100100010;
rgb[5814] = 24'b000110111011000000101001;
rgb[5815] = 24'b000111111100111000110000;
rgb[5816] = 24'b001100001101111101000001;
rgb[5817] = 24'b010011101110001101011100;
rgb[5818] = 24'b011010111110100001110111;
rgb[5819] = 24'b100010011110110010010010;
rgb[5820] = 24'b101001101111000110101101;
rgb[5821] = 24'b110001001111010111001000;
rgb[5822] = 24'b111000011111101011100011;
rgb[5823] = 24'b111111111111111111111111;
rgb[5824] = 24'b000000000000000000000000;
rgb[5825] = 24'b000000110001111000000101;
rgb[5826] = 24'b000001100011110100001011;
rgb[5827] = 24'b000010100101101100010001;
rgb[5828] = 24'b000011010111101000010111;
rgb[5829] = 24'b000100001001100100011101;
rgb[5830] = 24'b000101001011011100100011;
rgb[5831] = 24'b000101111101011000101001;
rgb[5832] = 24'b001010001110011100111010;
rgb[5833] = 24'b010001111110101001010110;
rgb[5834] = 24'b011001011110111001110010;
rgb[5835] = 24'b100001001111000110001110;
rgb[5836] = 24'b101000111111010010101010;
rgb[5837] = 24'b110000011111100011000110;
rgb[5838] = 24'b111000001111101111100010;
rgb[5839] = 24'b111111111111111111111111;
rgb[5840] = 24'b000000000000000000000000;
rgb[5841] = 24'b000000100001111100000101;
rgb[5842] = 24'b000001000011111100001010;
rgb[5843] = 24'b000001100101111100001111;
rgb[5844] = 24'b000010010111111000010100;
rgb[5845] = 24'b000010111001111000011001;
rgb[5846] = 24'b000011011011111000011110;
rgb[5847] = 24'b000011111101111000100011;
rgb[5848] = 24'b001000001110111100110100;
rgb[5849] = 24'b010000001111000101010001;
rgb[5850] = 24'b011000001111001101101110;
rgb[5851] = 24'b100000001111010110001011;
rgb[5852] = 24'b100111111111100010101000;
rgb[5853] = 24'b101111111111101011000101;
rgb[5854] = 24'b110111111111110011100010;
rgb[5855] = 24'b111111111111111111111111;
rgb[5856] = 24'b000000000000000000000000;
rgb[5857] = 24'b000000010010000000000100;
rgb[5858] = 24'b000000100100000100001000;
rgb[5859] = 24'b000000110110001000001100;
rgb[5860] = 24'b000001001000001100010000;
rgb[5861] = 24'b000001011010010000010100;
rgb[5862] = 24'b000001101100010100011000;
rgb[5863] = 24'b000001111110011000011101;
rgb[5864] = 24'b000110001111011100101110;
rgb[5865] = 24'b001110011111100001001011;
rgb[5866] = 24'b010110101111100101101001;
rgb[5867] = 24'b011110111111101010000111;
rgb[5868] = 24'b100111001111101110100101;
rgb[5869] = 24'b101111011111110011000011;
rgb[5870] = 24'b110111101111110111100001;
rgb[5871] = 24'b111111111111111111111111;
rgb[5872] = 24'b000000000000000000000000;
rgb[5873] = 24'b000000000010001000000011;
rgb[5874] = 24'b000000000100010000000110;
rgb[5875] = 24'b000000000110011000001001;
rgb[5876] = 24'b000000001000100000001100;
rgb[5877] = 24'b000000001010101000010000;
rgb[5878] = 24'b000000001100110000010011;
rgb[5879] = 24'b000000001110111000010110;
rgb[5880] = 24'b000100011111111000100111;
rgb[5881] = 24'b001100101111111101000110;
rgb[5882] = 24'b010101011111111001100101;
rgb[5883] = 24'b011101101111111110000011;
rgb[5884] = 24'b100110011111111110100010;
rgb[5885] = 24'b101110111111111111000001;
rgb[5886] = 24'b110111011111111111100000;
rgb[5887] = 24'b111111111111111111111111;
rgb[5888] = 24'b000000000000000000000000;
rgb[5889] = 24'b000100010001000100010001;
rgb[5890] = 24'b001000100010001000100010;
rgb[5891] = 24'b001100110011001100110011;
rgb[5892] = 24'b010001000100010001000100;
rgb[5893] = 24'b010101010101010101010101;
rgb[5894] = 24'b011001100110011001100110;
rgb[5895] = 24'b011101110111011101110111;
rgb[5896] = 24'b100010001000100010001000;
rgb[5897] = 24'b100110011001100110011001;
rgb[5898] = 24'b101010101010101010101010;
rgb[5899] = 24'b101110111011101110111011;
rgb[5900] = 24'b110011001100110011001100;
rgb[5901] = 24'b110111011101110111011101;
rgb[5902] = 24'b111011101110111011101110;
rgb[5903] = 24'b111111111111111111111111;
rgb[5904] = 24'b000000000000000000000000;
rgb[5905] = 24'b000011110001001000010000;
rgb[5906] = 24'b000111110010010000100000;
rgb[5907] = 24'b001011110011011000110000;
rgb[5908] = 24'b001111110100100001000001;
rgb[5909] = 24'b010011110101101001010001;
rgb[5910] = 24'b010111110110110001100001;
rgb[5911] = 24'b011011110111111001110010;
rgb[5912] = 24'b100000001000111110000011;
rgb[5913] = 24'b100100101001111110010100;
rgb[5914] = 24'b101001001010111110100110;
rgb[5915] = 24'b101101101011111110111000;
rgb[5916] = 24'b110010001100111111001001;
rgb[5917] = 24'b110110101101111111011011;
rgb[5918] = 24'b111011001110111111101101;
rgb[5919] = 24'b111111111111111111111111;
rgb[5920] = 24'b000000000000000000000000;
rgb[5921] = 24'b000011100001001100001111;
rgb[5922] = 24'b000111010010011000011111;
rgb[5923] = 24'b001011000011100100101110;
rgb[5924] = 24'b001110100100110100111110;
rgb[5925] = 24'b010010010110000001001101;
rgb[5926] = 24'b010110000111001101011101;
rgb[5927] = 24'b011001111000011001101101;
rgb[5928] = 24'b011110001001011101111110;
rgb[5929] = 24'b100010111010011010010000;
rgb[5930] = 24'b100111101011010110100010;
rgb[5931] = 24'b101100011100010010110101;
rgb[5932] = 24'b110001011101001011000111;
rgb[5933] = 24'b110110001110000111011010;
rgb[5934] = 24'b111010111111000011101100;
rgb[5935] = 24'b111111111111111111111111;
rgb[5936] = 24'b000000000000000000000000;
rgb[5937] = 24'b000011010001010000001110;
rgb[5938] = 24'b000110110010100000011101;
rgb[5939] = 24'b001010000011110100101100;
rgb[5940] = 24'b001101100101000100111011;
rgb[5941] = 24'b010001000110010101001010;
rgb[5942] = 24'b010100010111101001011001;
rgb[5943] = 24'b010111111000111001101000;
rgb[5944] = 24'b011100001001111101111001;
rgb[5945] = 24'b100001001010110110001100;
rgb[5946] = 24'b100110001011101110011111;
rgb[5947] = 24'b101011011100100010110010;
rgb[5948] = 24'b110000011101011011000101;
rgb[5949] = 24'b110101101110001111011000;
rgb[5950] = 24'b111010101111000111101011;
rgb[5951] = 24'b111111111111111111111111;
rgb[5952] = 24'b000000000000000000000000;
rgb[5953] = 24'b000011000001010100001110;
rgb[5954] = 24'b000110000010101100011100;
rgb[5955] = 24'b001001010100000000101010;
rgb[5956] = 24'b001100010101011000111000;
rgb[5957] = 24'b001111100110101101000110;
rgb[5958] = 24'b010010101000000101010101;
rgb[5959] = 24'b010101111001011001100011;
rgb[5960] = 24'b011010001010011101110100;
rgb[5961] = 24'b011111011011010010001000;
rgb[5962] = 24'b100100111100000010011011;
rgb[5963] = 24'b101010001100110110101111;
rgb[5964] = 24'b101111101101100111000011;
rgb[5965] = 24'b110100111110011011010111;
rgb[5966] = 24'b111010011111001011101011;
rgb[5967] = 24'b111111111111111111111111;
rgb[5968] = 24'b000000000000000000000000;
rgb[5969] = 24'b000010110001011000001101;
rgb[5970] = 24'b000101100010110100011010;
rgb[5971] = 24'b001000100100010000101000;
rgb[5972] = 24'b001011010101101000110101;
rgb[5973] = 24'b001110000111000101000011;
rgb[5974] = 24'b010001001000100001010000;
rgb[5975] = 24'b010011111001111001011110;
rgb[5976] = 24'b011000001010111101101111;
rgb[5977] = 24'b011101101011101110000011;
rgb[5978] = 24'b100011011100011010011000;
rgb[5979] = 24'b101001001101000110101100;
rgb[5980] = 24'b101110111101110111000001;
rgb[5981] = 24'b110100011110100011010101;
rgb[5982] = 24'b111010001111001111101010;
rgb[5983] = 24'b111111111111111111111111;
rgb[5984] = 24'b000000000000000000000000;
rgb[5985] = 24'b000010100001011100001100;
rgb[5986] = 24'b000101000010111100011001;
rgb[5987] = 24'b000111100100011100100110;
rgb[5988] = 24'b001010000101111100110011;
rgb[5989] = 24'b001100110111011000111111;
rgb[5990] = 24'b001111011000111001001100;
rgb[5991] = 24'b010001111010011001011001;
rgb[5992] = 24'b010110001011011101101010;
rgb[5993] = 24'b011100001100000101111111;
rgb[5994] = 24'b100001111100110010010100;
rgb[5995] = 24'b100111111101011010101010;
rgb[5996] = 24'b101101111110000010111111;
rgb[5997] = 24'b110011111110101011010100;
rgb[5998] = 24'b111001111111010011101001;
rgb[5999] = 24'b111111111111111011111111;
rgb[6000] = 24'b000000000000000000000000;
rgb[6001] = 24'b000010010001100000001100;
rgb[6002] = 24'b000100100011000100011000;
rgb[6003] = 24'b000110110100101000100100;
rgb[6004] = 24'b001001000110001100110000;
rgb[6005] = 24'b001011010111110000111100;
rgb[6006] = 24'b001101101001010101001000;
rgb[6007] = 24'b001111111010111001010100;
rgb[6008] = 24'b010100001011111101100101;
rgb[6009] = 24'b011010011100100001111011;
rgb[6010] = 24'b100000101101000110010001;
rgb[6011] = 24'b100110111101101010100111;
rgb[6012] = 24'b101101001110001110111101;
rgb[6013] = 24'b110011011110110011010011;
rgb[6014] = 24'b111001101111010111101001;
rgb[6015] = 24'b111111111111111111111111;
rgb[6016] = 24'b000000000000000000000000;
rgb[6017] = 24'b000001110001101000001011;
rgb[6018] = 24'b000011110011010000010110;
rgb[6019] = 24'b000101110100111000100010;
rgb[6020] = 24'b000111110110100000101101;
rgb[6021] = 24'b001001111000001000111000;
rgb[6022] = 24'b001011111001110001000100;
rgb[6023] = 24'b001101111011011001001111;
rgb[6024] = 24'b010010001100011101100000;
rgb[6025] = 24'b011000101100111101110111;
rgb[6026] = 24'b011111001101011110001101;
rgb[6027] = 24'b100101101101111110100100;
rgb[6028] = 24'b101100001110011110111011;
rgb[6029] = 24'b110010101110111111010001;
rgb[6030] = 24'b111001001111011111101000;
rgb[6031] = 24'b111111111111111011111111;
rgb[6032] = 24'b000000000000000000000000;
rgb[6033] = 24'b000001100001101100001010;
rgb[6034] = 24'b000011010011011000010101;
rgb[6035] = 24'b000101000101000100100000;
rgb[6036] = 24'b000110110110110000101010;
rgb[6037] = 24'b001000011000100000110101;
rgb[6038] = 24'b001010001010001101000000;
rgb[6039] = 24'b001011111011111001001010;
rgb[6040] = 24'b010000001100111101011011;
rgb[6041] = 24'b010110111101011001110011;
rgb[6042] = 24'b011101101101110110001010;
rgb[6043] = 24'b100100101110001110100001;
rgb[6044] = 24'b101011011110101010111001;
rgb[6045] = 24'b110010001111000111010000;
rgb[6046] = 24'b111000111111100011100111;
rgb[6047] = 24'b111111111111111111111111;
rgb[6048] = 24'b000000000000000000000000;
rgb[6049] = 24'b000001010001110000001001;
rgb[6050] = 24'b000010110011100000010011;
rgb[6051] = 24'b000100010101010100011101;
rgb[6052] = 24'b000101100111000100100111;
rgb[6053] = 24'b000111001000110100110001;
rgb[6054] = 24'b001000101010101000111011;
rgb[6055] = 24'b001001111100011001000101;
rgb[6056] = 24'b001110001101011101010110;
rgb[6057] = 24'b010101001101110101101110;
rgb[6058] = 24'b011100011110001010000110;
rgb[6059] = 24'b100011011110100010011110;
rgb[6060] = 24'b101010101110111010110110;
rgb[6061] = 24'b110001101111001111001110;
rgb[6062] = 24'b111000101111100111100110;
rgb[6063] = 24'b111111111111111011111111;
rgb[6064] = 24'b000000000000000000000000;
rgb[6065] = 24'b000001000001110100001001;
rgb[6066] = 24'b000010010011101000010010;
rgb[6067] = 24'b000011010101100000011011;
rgb[6068] = 24'b000100100111010100100101;
rgb[6069] = 24'b000101101001001100101110;
rgb[6070] = 24'b000110111011000000110111;
rgb[6071] = 24'b000111111100111001000000;
rgb[6072] = 24'b001100001101111101010001;
rgb[6073] = 24'b010011101110001101101010;
rgb[6074] = 24'b011010111110100010000011;
rgb[6075] = 24'b100010011110110010011100;
rgb[6076] = 24'b101001101111000110110100;
rgb[6077] = 24'b110001001111010111001101;
rgb[6078] = 24'b111000011111101011100110;
rgb[6079] = 24'b111111111111111111111111;
rgb[6080] = 24'b000000000000000000000000;
rgb[6081] = 24'b000000110001111000001000;
rgb[6082] = 24'b000001100011110100010001;
rgb[6083] = 24'b000010100101101100011001;
rgb[6084] = 24'b000011010111101000100010;
rgb[6085] = 24'b000100001001100100101010;
rgb[6086] = 24'b000101001011011100110011;
rgb[6087] = 24'b000101111101011000111100;
rgb[6088] = 24'b001010001110011101001101;
rgb[6089] = 24'b010001111110101001100110;
rgb[6090] = 24'b011001011110111001111111;
rgb[6091] = 24'b100001001111000110011001;
rgb[6092] = 24'b101000111111010010110010;
rgb[6093] = 24'b110000011111100011001100;
rgb[6094] = 24'b111000001111101111100101;
rgb[6095] = 24'b111111111111111111111111;
rgb[6096] = 24'b000000000000000000000000;
rgb[6097] = 24'b000000100001111100000111;
rgb[6098] = 24'b000001000011111100001111;
rgb[6099] = 24'b000001100101111100010111;
rgb[6100] = 24'b000010010111111000011111;
rgb[6101] = 24'b000010111001111000100111;
rgb[6102] = 24'b000011011011111000101111;
rgb[6103] = 24'b000011111101111000110111;
rgb[6104] = 24'b001000001110111101001000;
rgb[6105] = 24'b010000001111000101100010;
rgb[6106] = 24'b011000001111001101111100;
rgb[6107] = 24'b100000001111010110010110;
rgb[6108] = 24'b100111111111100010110000;
rgb[6109] = 24'b101111111111101011001010;
rgb[6110] = 24'b110111111111110011100100;
rgb[6111] = 24'b111111111111111111111111;
rgb[6112] = 24'b000000000000000000000000;
rgb[6113] = 24'b000000010010000000000111;
rgb[6114] = 24'b000000100100000100001110;
rgb[6115] = 24'b000000110110001000010101;
rgb[6116] = 24'b000001001000001100011100;
rgb[6117] = 24'b000001011010010000100011;
rgb[6118] = 24'b000001101100010100101011;
rgb[6119] = 24'b000001111110011000110010;
rgb[6120] = 24'b000110001111011101000011;
rgb[6121] = 24'b001110011111100001011110;
rgb[6122] = 24'b010110101111100101111000;
rgb[6123] = 24'b011110111111101010010011;
rgb[6124] = 24'b100111001111101110101110;
rgb[6125] = 24'b101111011111110011001001;
rgb[6126] = 24'b110111101111110111100100;
rgb[6127] = 24'b111111111111111111111111;
rgb[6128] = 24'b000000000000000000000000;
rgb[6129] = 24'b000000000010001000000110;
rgb[6130] = 24'b000000000100010000001100;
rgb[6131] = 24'b000000000110011000010011;
rgb[6132] = 24'b000000001000100000011001;
rgb[6133] = 24'b000000001010101000100000;
rgb[6134] = 24'b000000001100110000100110;
rgb[6135] = 24'b000000001110111000101101;
rgb[6136] = 24'b000100011111111000111110;
rgb[6137] = 24'b001100101111111101011001;
rgb[6138] = 24'b010101011111111001110101;
rgb[6139] = 24'b011101101111111110010000;
rgb[6140] = 24'b100110011111111110101100;
rgb[6141] = 24'b101110111111111111000111;
rgb[6142] = 24'b110111011111111111100011;
rgb[6143] = 24'b111111111111111111111111;
rgb[6144] = 24'b000000000000000000000000;
rgb[6145] = 24'b000100010001000100010001;
rgb[6146] = 24'b001000100010001000100010;
rgb[6147] = 24'b001100110011001100110011;
rgb[6148] = 24'b010001000100010001000100;
rgb[6149] = 24'b010101010101010101010101;
rgb[6150] = 24'b011001100110011001100110;
rgb[6151] = 24'b011101110111011101110111;
rgb[6152] = 24'b100010001000100010001000;
rgb[6153] = 24'b100110011001100110011001;
rgb[6154] = 24'b101010101010101010101010;
rgb[6155] = 24'b101110111011101110111011;
rgb[6156] = 24'b110011001100110011001100;
rgb[6157] = 24'b110111011101110111011101;
rgb[6158] = 24'b111011101110111011101110;
rgb[6159] = 24'b111111111111111111111111;
rgb[6160] = 24'b000000000000000000000000;
rgb[6161] = 24'b000011110001001000010000;
rgb[6162] = 24'b000111110010010000100001;
rgb[6163] = 24'b001011110011011000110001;
rgb[6164] = 24'b001111110100100001000010;
rgb[6165] = 24'b010011110101101001010010;
rgb[6166] = 24'b010111110110110001100011;
rgb[6167] = 24'b011011110111111001110011;
rgb[6168] = 24'b100000001000111110000100;
rgb[6169] = 24'b100100101001111110010110;
rgb[6170] = 24'b101001001010111110100111;
rgb[6171] = 24'b101101101011111110111001;
rgb[6172] = 24'b110010001100111111001010;
rgb[6173] = 24'b110110101101111111011100;
rgb[6174] = 24'b111011001110111111101101;
rgb[6175] = 24'b111111111111111111111111;
rgb[6176] = 24'b000000000000000000000000;
rgb[6177] = 24'b000011100001001100010000;
rgb[6178] = 24'b000111010010011000100000;
rgb[6179] = 24'b001011000011100100110000;
rgb[6180] = 24'b001110100100110101000000;
rgb[6181] = 24'b010010010110000001010000;
rgb[6182] = 24'b010110000111001101100000;
rgb[6183] = 24'b011001111000011001110000;
rgb[6184] = 24'b011110001001011110000001;
rgb[6185] = 24'b100010111010011010010011;
rgb[6186] = 24'b100111101011010110100101;
rgb[6187] = 24'b101100011100010010110111;
rgb[6188] = 24'b110001011101001011001001;
rgb[6189] = 24'b110110001110000111011011;
rgb[6190] = 24'b111010111111000011101101;
rgb[6191] = 24'b111111111111111111111111;
rgb[6192] = 24'b000000000000000000000000;
rgb[6193] = 24'b000011010001010000001111;
rgb[6194] = 24'b000110110010100000011111;
rgb[6195] = 24'b001010000011110100101110;
rgb[6196] = 24'b001101100101000100111110;
rgb[6197] = 24'b010001000110010101001101;
rgb[6198] = 24'b010100010111101001011101;
rgb[6199] = 24'b010111111000111001101100;
rgb[6200] = 24'b011100001001111101111101;
rgb[6201] = 24'b100001001010110110010000;
rgb[6202] = 24'b100110001011101110100010;
rgb[6203] = 24'b101011011100100010110101;
rgb[6204] = 24'b110000011101011011000111;
rgb[6205] = 24'b110101101110001111011010;
rgb[6206] = 24'b111010101111000111101100;
rgb[6207] = 24'b111111111111111111111111;
rgb[6208] = 24'b000000000000000000000000;
rgb[6209] = 24'b000011000001010100001111;
rgb[6210] = 24'b000110000010101100011110;
rgb[6211] = 24'b001001010100000000101101;
rgb[6212] = 24'b001100010101011000111100;
rgb[6213] = 24'b001111100110101101001011;
rgb[6214] = 24'b010010101000000101011010;
rgb[6215] = 24'b010101111001011001101001;
rgb[6216] = 24'b011010001010011101111010;
rgb[6217] = 24'b011111011011010010001101;
rgb[6218] = 24'b100100111100000010100000;
rgb[6219] = 24'b101010001100110110110011;
rgb[6220] = 24'b101111101101100111000110;
rgb[6221] = 24'b110100111110011011011001;
rgb[6222] = 24'b111010011111001011101100;
rgb[6223] = 24'b111111111111111111111111;
rgb[6224] = 24'b000000000000000000000000;
rgb[6225] = 24'b000010110001011000001110;
rgb[6226] = 24'b000101100010110100011101;
rgb[6227] = 24'b001000100100010000101011;
rgb[6228] = 24'b001011010101101000111010;
rgb[6229] = 24'b001110000111000101001000;
rgb[6230] = 24'b010001001000100001010111;
rgb[6231] = 24'b010011111001111001100110;
rgb[6232] = 24'b011000001010111101110111;
rgb[6233] = 24'b011101101011101110001010;
rgb[6234] = 24'b100011011100011010011101;
rgb[6235] = 24'b101001001101000110110001;
rgb[6236] = 24'b101110111101110111000100;
rgb[6237] = 24'b110100011110100011011000;
rgb[6238] = 24'b111010001111001111101011;
rgb[6239] = 24'b111111111111111111111111;
rgb[6240] = 24'b000000000000000000000000;
rgb[6241] = 24'b000010100001011100001110;
rgb[6242] = 24'b000101000010111100011100;
rgb[6243] = 24'b000111100100011100101010;
rgb[6244] = 24'b001010000101111100111000;
rgb[6245] = 24'b001100110111011001000110;
rgb[6246] = 24'b001111011000111001010100;
rgb[6247] = 24'b010001111010011001100010;
rgb[6248] = 24'b010110001011011101110011;
rgb[6249] = 24'b011100001100000110000111;
rgb[6250] = 24'b100001111100110010011011;
rgb[6251] = 24'b100111111101011010101111;
rgb[6252] = 24'b101101111110000011000011;
rgb[6253] = 24'b110011111110101011010111;
rgb[6254] = 24'b111001111111010011101011;
rgb[6255] = 24'b111111111111111011111111;
rgb[6256] = 24'b000000000000000000000000;
rgb[6257] = 24'b000010010001100000001101;
rgb[6258] = 24'b000100100011000100011011;
rgb[6259] = 24'b000110110100101000101000;
rgb[6260] = 24'b001001000110001100110110;
rgb[6261] = 24'b001011010111110001000011;
rgb[6262] = 24'b001101101001010101010001;
rgb[6263] = 24'b001111111010111001011111;
rgb[6264] = 24'b010100001011111101110000;
rgb[6265] = 24'b011010011100100010000100;
rgb[6266] = 24'b100000101101000110011001;
rgb[6267] = 24'b100110111101101010101101;
rgb[6268] = 24'b101101001110001111000001;
rgb[6269] = 24'b110011011110110011010110;
rgb[6270] = 24'b111001101111010111101010;
rgb[6271] = 24'b111111111111111111111111;
rgb[6272] = 24'b000000000000000000000000;
rgb[6273] = 24'b000001110001101000001101;
rgb[6274] = 24'b000011110011010000011010;
rgb[6275] = 24'b000101110100111000100111;
rgb[6276] = 24'b000111110110100000110100;
rgb[6277] = 24'b001001111000001001000001;
rgb[6278] = 24'b001011111001110001001110;
rgb[6279] = 24'b001101111011011001011011;
rgb[6280] = 24'b010010001100011101101100;
rgb[6281] = 24'b011000101100111110000001;
rgb[6282] = 24'b011111001101011110010110;
rgb[6283] = 24'b100101101101111110101011;
rgb[6284] = 24'b101100001110011111000000;
rgb[6285] = 24'b110010101110111111010101;
rgb[6286] = 24'b111001001111011111101010;
rgb[6287] = 24'b111111111111111011111111;
rgb[6288] = 24'b000000000000000000000000;
rgb[6289] = 24'b000001100001101100001100;
rgb[6290] = 24'b000011010011011000011001;
rgb[6291] = 24'b000101000101000100100101;
rgb[6292] = 24'b000110110110110000110010;
rgb[6293] = 24'b001000011000100000111111;
rgb[6294] = 24'b001010001010001101001011;
rgb[6295] = 24'b001011111011111001011000;
rgb[6296] = 24'b010000001100111101101001;
rgb[6297] = 24'b010110111101011001111110;
rgb[6298] = 24'b011101101101110110010100;
rgb[6299] = 24'b100100101110001110101001;
rgb[6300] = 24'b101011011110101010111110;
rgb[6301] = 24'b110010001111000111010100;
rgb[6302] = 24'b111000111111100011101001;
rgb[6303] = 24'b111111111111111111111111;
rgb[6304] = 24'b000000000000000000000000;
rgb[6305] = 24'b000001010001110000001100;
rgb[6306] = 24'b000010110011100000011000;
rgb[6307] = 24'b000100010101010100100100;
rgb[6308] = 24'b000101100111000100110000;
rgb[6309] = 24'b000111001000110100111100;
rgb[6310] = 24'b001000101010101001001000;
rgb[6311] = 24'b001001111100011001010101;
rgb[6312] = 24'b001110001101011101100101;
rgb[6313] = 24'b010101001101110101111011;
rgb[6314] = 24'b011100011110001010010001;
rgb[6315] = 24'b100011011110100010100111;
rgb[6316] = 24'b101010101110111010111101;
rgb[6317] = 24'b110001101111001111010011;
rgb[6318] = 24'b111000101111100111101001;
rgb[6319] = 24'b111111111111111011111111;
rgb[6320] = 24'b000000000000000000000000;
rgb[6321] = 24'b000001000001110100001011;
rgb[6322] = 24'b000010010011101000010111;
rgb[6323] = 24'b000011010101100000100010;
rgb[6324] = 24'b000100100111010100101110;
rgb[6325] = 24'b000101101001001100111010;
rgb[6326] = 24'b000110111011000001000101;
rgb[6327] = 24'b000111111100111001010001;
rgb[6328] = 24'b001100001101111101100010;
rgb[6329] = 24'b010011101110001101111000;
rgb[6330] = 24'b011010111110100010001111;
rgb[6331] = 24'b100010011110110010100101;
rgb[6332] = 24'b101001101111000110111011;
rgb[6333] = 24'b110001001111010111010010;
rgb[6334] = 24'b111000011111101011101000;
rgb[6335] = 24'b111111111111111111111111;
rgb[6336] = 24'b000000000000000000000000;
rgb[6337] = 24'b000000110001111000001011;
rgb[6338] = 24'b000001100011110100010110;
rgb[6339] = 24'b000010100101101100100001;
rgb[6340] = 24'b000011010111101000101100;
rgb[6341] = 24'b000100001001100100110111;
rgb[6342] = 24'b000101001011011101000011;
rgb[6343] = 24'b000101111101011001001110;
rgb[6344] = 24'b001010001110011101011111;
rgb[6345] = 24'b010001111110101001110110;
rgb[6346] = 24'b011001011110111010001100;
rgb[6347] = 24'b100001001111000110100011;
rgb[6348] = 24'b101000111111010010111010;
rgb[6349] = 24'b110000011111100011010001;
rgb[6350] = 24'b111000001111101111101000;
rgb[6351] = 24'b111111111111111111111111;
rgb[6352] = 24'b000000000000000000000000;
rgb[6353] = 24'b000000100001111100001010;
rgb[6354] = 24'b000001000011111100010101;
rgb[6355] = 24'b000001100101111100100000;
rgb[6356] = 24'b000010010111111000101010;
rgb[6357] = 24'b000010111001111000110101;
rgb[6358] = 24'b000011011011111001000000;
rgb[6359] = 24'b000011111101111001001010;
rgb[6360] = 24'b001000001110111101011011;
rgb[6361] = 24'b010000001111000101110011;
rgb[6362] = 24'b011000001111001110001010;
rgb[6363] = 24'b100000001111010110100001;
rgb[6364] = 24'b100111111111100010111001;
rgb[6365] = 24'b101111111111101011010000;
rgb[6366] = 24'b110111111111110011100111;
rgb[6367] = 24'b111111111111111111111111;
rgb[6368] = 24'b000000000000000000000000;
rgb[6369] = 24'b000000010010000000001010;
rgb[6370] = 24'b000000100100000100010100;
rgb[6371] = 24'b000000110110001000011110;
rgb[6372] = 24'b000001001000001100101000;
rgb[6373] = 24'b000001011010010000110011;
rgb[6374] = 24'b000001101100010100111101;
rgb[6375] = 24'b000001111110011001000111;
rgb[6376] = 24'b000110001111011101011000;
rgb[6377] = 24'b001110011111100001110000;
rgb[6378] = 24'b010110101111100110000111;
rgb[6379] = 24'b011110111111101010011111;
rgb[6380] = 24'b100111001111101110110111;
rgb[6381] = 24'b101111011111110011001111;
rgb[6382] = 24'b110111101111110111100111;
rgb[6383] = 24'b111111111111111111111111;
rgb[6384] = 24'b000000000000000000000000;
rgb[6385] = 24'b000000000010001000001001;
rgb[6386] = 24'b000000000100010000010011;
rgb[6387] = 24'b000000000110011000011101;
rgb[6388] = 24'b000000001000100000100110;
rgb[6389] = 24'b000000001010101000110000;
rgb[6390] = 24'b000000001100110000111010;
rgb[6391] = 24'b000000001110111001000100;
rgb[6392] = 24'b000100011111111001010101;
rgb[6393] = 24'b001100101111111101101101;
rgb[6394] = 24'b010101011111111010000101;
rgb[6395] = 24'b011101101111111110011101;
rgb[6396] = 24'b100110011111111110110110;
rgb[6397] = 24'b101110111111111111001110;
rgb[6398] = 24'b110111011111111111100110;
rgb[6399] = 24'b111111111111111111111111;
rgb[6400] = 24'b000000000000000000000000;
rgb[6401] = 24'b000100010001000100010001;
rgb[6402] = 24'b001000100010001000100010;
rgb[6403] = 24'b001100110011001100110011;
rgb[6404] = 24'b010001000100010001000100;
rgb[6405] = 24'b010101010101010101010101;
rgb[6406] = 24'b011001100110011001100110;
rgb[6407] = 24'b011101110111011101110111;
rgb[6408] = 24'b100010001000100010001000;
rgb[6409] = 24'b100110011001100110011001;
rgb[6410] = 24'b101010101010101010101010;
rgb[6411] = 24'b101110111011101110111011;
rgb[6412] = 24'b110011001100110011001100;
rgb[6413] = 24'b110111011101110111011101;
rgb[6414] = 24'b111011101110111011101110;
rgb[6415] = 24'b111111111111111111111111;
rgb[6416] = 24'b000000000000000000000000;
rgb[6417] = 24'b000011110001001000010000;
rgb[6418] = 24'b000111110010010000100001;
rgb[6419] = 24'b001011110011011000110010;
rgb[6420] = 24'b001111110100100001000010;
rgb[6421] = 24'b010011110101101001010011;
rgb[6422] = 24'b010111110110110001100100;
rgb[6423] = 24'b011011110111111001110101;
rgb[6424] = 24'b100000001000111110000110;
rgb[6425] = 24'b100100101001111110010111;
rgb[6426] = 24'b101001001010111110101000;
rgb[6427] = 24'b101101101011111110111001;
rgb[6428] = 24'b110010001100111111001011;
rgb[6429] = 24'b110110101101111111011100;
rgb[6430] = 24'b111011001110111111101101;
rgb[6431] = 24'b111111111111111111111111;
rgb[6432] = 24'b000000000000000000000000;
rgb[6433] = 24'b000011100001001100010000;
rgb[6434] = 24'b000111010010011000100000;
rgb[6435] = 24'b001011000011100100110001;
rgb[6436] = 24'b001110100100110101000001;
rgb[6437] = 24'b010010010110000001010010;
rgb[6438] = 24'b010110000111001101100010;
rgb[6439] = 24'b011001111000011001110011;
rgb[6440] = 24'b011110001001011110000100;
rgb[6441] = 24'b100010111010011010010101;
rgb[6442] = 24'b100111101011010110100111;
rgb[6443] = 24'b101100011100010010111000;
rgb[6444] = 24'b110001011101001011001010;
rgb[6445] = 24'b110110001110000111011011;
rgb[6446] = 24'b111010111111000011101101;
rgb[6447] = 24'b111111111111111111111111;
rgb[6448] = 24'b000000000000000000000000;
rgb[6449] = 24'b000011010001010000010000;
rgb[6450] = 24'b000110110010100000100000;
rgb[6451] = 24'b001010000011110100110000;
rgb[6452] = 24'b001101100101000101000000;
rgb[6453] = 24'b010001000110010101010000;
rgb[6454] = 24'b010100010111101001100001;
rgb[6455] = 24'b010111111000111001110001;
rgb[6456] = 24'b011100001001111110000010;
rgb[6457] = 24'b100001001010110110010100;
rgb[6458] = 24'b100110001011101110100101;
rgb[6459] = 24'b101011011100100010110111;
rgb[6460] = 24'b110000011101011011001001;
rgb[6461] = 24'b110101101110001111011011;
rgb[6462] = 24'b111010101111000111101101;
rgb[6463] = 24'b111111111111111111111111;
rgb[6464] = 24'b000000000000000000000000;
rgb[6465] = 24'b000011000001010100001111;
rgb[6466] = 24'b000110000010101100011111;
rgb[6467] = 24'b001001010100000000101111;
rgb[6468] = 24'b001100010101011000111111;
rgb[6469] = 24'b001111100110101101001111;
rgb[6470] = 24'b010010101000000101011111;
rgb[6471] = 24'b010101111001011001101111;
rgb[6472] = 24'b011010001010011110000000;
rgb[6473] = 24'b011111011011010010010010;
rgb[6474] = 24'b100100111100000010100100;
rgb[6475] = 24'b101010001100110110110110;
rgb[6476] = 24'b101111101101100111001000;
rgb[6477] = 24'b110100111110011011011010;
rgb[6478] = 24'b111010011111001011101100;
rgb[6479] = 24'b111111111111111111111111;
rgb[6480] = 24'b000000000000000000000000;
rgb[6481] = 24'b000010110001011000001111;
rgb[6482] = 24'b000101100010110100011111;
rgb[6483] = 24'b001000100100010000101110;
rgb[6484] = 24'b001011010101101000111110;
rgb[6485] = 24'b001110000111000101001110;
rgb[6486] = 24'b010001001000100001011101;
rgb[6487] = 24'b010011111001111001101101;
rgb[6488] = 24'b011000001010111101111110;
rgb[6489] = 24'b011101101011101110010000;
rgb[6490] = 24'b100011011100011010100011;
rgb[6491] = 24'b101001001101000110110101;
rgb[6492] = 24'b101110111101110111000111;
rgb[6493] = 24'b110100011110100011011010;
rgb[6494] = 24'b111010001111001111101100;
rgb[6495] = 24'b111111111111111111111111;
rgb[6496] = 24'b000000000000000000000000;
rgb[6497] = 24'b000010100001011100001111;
rgb[6498] = 24'b000101000010111100011110;
rgb[6499] = 24'b000111100100011100101110;
rgb[6500] = 24'b001010000101111100111101;
rgb[6501] = 24'b001100110111011001001100;
rgb[6502] = 24'b001111011000111001011100;
rgb[6503] = 24'b010001111010011001101011;
rgb[6504] = 24'b010110001011011101111100;
rgb[6505] = 24'b011100001100000110001111;
rgb[6506] = 24'b100001111100110010100001;
rgb[6507] = 24'b100111111101011010110100;
rgb[6508] = 24'b101101111110000011000111;
rgb[6509] = 24'b110011111110101011011001;
rgb[6510] = 24'b111001111111010011101100;
rgb[6511] = 24'b111111111111111011111111;
rgb[6512] = 24'b000000000000000000000000;
rgb[6513] = 24'b000010010001100000001111;
rgb[6514] = 24'b000100100011000100011110;
rgb[6515] = 24'b000110110100101000101101;
rgb[6516] = 24'b001001000110001100111100;
rgb[6517] = 24'b001011010111110001001011;
rgb[6518] = 24'b001101101001010101011010;
rgb[6519] = 24'b001111111010111001101001;
rgb[6520] = 24'b010100001011111101111010;
rgb[6521] = 24'b011010011100100010001101;
rgb[6522] = 24'b100000101101000110100000;
rgb[6523] = 24'b100110111101101010110011;
rgb[6524] = 24'b101101001110001111000110;
rgb[6525] = 24'b110011011110110011011001;
rgb[6526] = 24'b111001101111010111101100;
rgb[6527] = 24'b111111111111111111111111;
rgb[6528] = 24'b000000000000000000000000;
rgb[6529] = 24'b000001110001101000001110;
rgb[6530] = 24'b000011110011010000011101;
rgb[6531] = 24'b000101110100111000101100;
rgb[6532] = 24'b000111110110100000111011;
rgb[6533] = 24'b001001111000001001001010;
rgb[6534] = 24'b001011111001110001011001;
rgb[6535] = 24'b001101111011011001100111;
rgb[6536] = 24'b010010001100011101111000;
rgb[6537] = 24'b011000101100111110001100;
rgb[6538] = 24'b011111001101011110011111;
rgb[6539] = 24'b100101101101111110110010;
rgb[6540] = 24'b101100001110011111000101;
rgb[6541] = 24'b110010101110111111011000;
rgb[6542] = 24'b111001001111011111101011;
rgb[6543] = 24'b111111111111111011111111;
rgb[6544] = 24'b000000000000000000000000;
rgb[6545] = 24'b000001100001101100001110;
rgb[6546] = 24'b000011010011011000011101;
rgb[6547] = 24'b000101000101000100101011;
rgb[6548] = 24'b000110110110110000111010;
rgb[6549] = 24'b001000011000100001001000;
rgb[6550] = 24'b001010001010001101010111;
rgb[6551] = 24'b001011111011111001100101;
rgb[6552] = 24'b010000001100111101110111;
rgb[6553] = 24'b010110111101011010001010;
rgb[6554] = 24'b011101101101110110011101;
rgb[6555] = 24'b100100101110001110110001;
rgb[6556] = 24'b101011011110101011000100;
rgb[6557] = 24'b110010001111000111011000;
rgb[6558] = 24'b111000111111100011101011;
rgb[6559] = 24'b111111111111111111111111;
rgb[6560] = 24'b000000000000000000000000;
rgb[6561] = 24'b000001010001110000001110;
rgb[6562] = 24'b000010110011100000011100;
rgb[6563] = 24'b000100010101010100101010;
rgb[6564] = 24'b000101100111000100111001;
rgb[6565] = 24'b000111001000110101000111;
rgb[6566] = 24'b001000101010101001010101;
rgb[6567] = 24'b001001111100011001100100;
rgb[6568] = 24'b001110001101011101110101;
rgb[6569] = 24'b010101001101110110001000;
rgb[6570] = 24'b011100011110001010011100;
rgb[6571] = 24'b100011011110100010110000;
rgb[6572] = 24'b101010101110111011000011;
rgb[6573] = 24'b110001101111001111010111;
rgb[6574] = 24'b111000101111100111101011;
rgb[6575] = 24'b111111111111111011111111;
rgb[6576] = 24'b000000000000000000000000;
rgb[6577] = 24'b000001000001110100001110;
rgb[6578] = 24'b000010010011101000011100;
rgb[6579] = 24'b000011010101100000101010;
rgb[6580] = 24'b000100100111010100111000;
rgb[6581] = 24'b000101101001001101000110;
rgb[6582] = 24'b000110111011000001010100;
rgb[6583] = 24'b000111111100111001100010;
rgb[6584] = 24'b001100001101111101110011;
rgb[6585] = 24'b010011101110001110000111;
rgb[6586] = 24'b011010111110100010011011;
rgb[6587] = 24'b100010011110110010101111;
rgb[6588] = 24'b101001101111000111000011;
rgb[6589] = 24'b110001001111010111010111;
rgb[6590] = 24'b111000011111101011101011;
rgb[6591] = 24'b111111111111111111111111;
rgb[6592] = 24'b000000000000000000000000;
rgb[6593] = 24'b000000110001111000001101;
rgb[6594] = 24'b000001100011110100011011;
rgb[6595] = 24'b000010100101101100101001;
rgb[6596] = 24'b000011010111101000110111;
rgb[6597] = 24'b000100001001100101000100;
rgb[6598] = 24'b000101001011011101010010;
rgb[6599] = 24'b000101111101011001100000;
rgb[6600] = 24'b001010001110011101110001;
rgb[6601] = 24'b010001111110101010000101;
rgb[6602] = 24'b011001011110111010011001;
rgb[6603] = 24'b100001001111000110101110;
rgb[6604] = 24'b101000111111010011000010;
rgb[6605] = 24'b110000011111100011010110;
rgb[6606] = 24'b111000001111101111101010;
rgb[6607] = 24'b111111111111111111111111;
rgb[6608] = 24'b000000000000000000000000;
rgb[6609] = 24'b000000100001111100001101;
rgb[6610] = 24'b000001000011111100011010;
rgb[6611] = 24'b000001100101111100101000;
rgb[6612] = 24'b000010010111111000110101;
rgb[6613] = 24'b000010111001111001000011;
rgb[6614] = 24'b000011011011111001010000;
rgb[6615] = 24'b000011111101111001011110;
rgb[6616] = 24'b001000001110111101101111;
rgb[6617] = 24'b010000001111000110000011;
rgb[6618] = 24'b011000001111001110011000;
rgb[6619] = 24'b100000001111010110101100;
rgb[6620] = 24'b100111111111100011000001;
rgb[6621] = 24'b101111111111101011010101;
rgb[6622] = 24'b110111111111110011101010;
rgb[6623] = 24'b111111111111111111111111;
rgb[6624] = 24'b000000000000000000000000;
rgb[6625] = 24'b000000010010000000001101;
rgb[6626] = 24'b000000100100000100011010;
rgb[6627] = 24'b000000110110001000100111;
rgb[6628] = 24'b000001001000001100110100;
rgb[6629] = 24'b000001011010010001000010;
rgb[6630] = 24'b000001101100010101001111;
rgb[6631] = 24'b000001111110011001011100;
rgb[6632] = 24'b000110001111011101101101;
rgb[6633] = 24'b001110011111100010000010;
rgb[6634] = 24'b010110101111100110010111;
rgb[6635] = 24'b011110111111101010101011;
rgb[6636] = 24'b100111001111101111000000;
rgb[6637] = 24'b101111011111110011010101;
rgb[6638] = 24'b110111101111110111101010;
rgb[6639] = 24'b111111111111111111111111;
rgb[6640] = 24'b000000000000000000000000;
rgb[6641] = 24'b000000000010001000001100;
rgb[6642] = 24'b000000000100010000011001;
rgb[6643] = 24'b000000000110011000100110;
rgb[6644] = 24'b000000001000100000110011;
rgb[6645] = 24'b000000001010101001000000;
rgb[6646] = 24'b000000001100110001001101;
rgb[6647] = 24'b000000001110111001011010;
rgb[6648] = 24'b000100011111111001101011;
rgb[6649] = 24'b001100101111111110000000;
rgb[6650] = 24'b010101011111111010010101;
rgb[6651] = 24'b011101101111111110101010;
rgb[6652] = 24'b100110011111111110111111;
rgb[6653] = 24'b101110111111111111010100;
rgb[6654] = 24'b110111011111111111101001;
rgb[6655] = 24'b111111111111111111111111;
rgb[6656] = 24'b000000000000000000000000;
rgb[6657] = 24'b000100010001000100010001;
rgb[6658] = 24'b001000100010001000100010;
rgb[6659] = 24'b001100110011001100110011;
rgb[6660] = 24'b010001000100010001000100;
rgb[6661] = 24'b010101010101010101010101;
rgb[6662] = 24'b011001100110011001100110;
rgb[6663] = 24'b011101110111011101110111;
rgb[6664] = 24'b100010001000100010001000;
rgb[6665] = 24'b100110011001100110011001;
rgb[6666] = 24'b101010101010101010101010;
rgb[6667] = 24'b101110111011101110111011;
rgb[6668] = 24'b110011001100110011001100;
rgb[6669] = 24'b110111011101110111011101;
rgb[6670] = 24'b111011101110111011101110;
rgb[6671] = 24'b111111111111111111111111;
rgb[6672] = 24'b000000000000000000000000;
rgb[6673] = 24'b000011110001001000010000;
rgb[6674] = 24'b000111110010010000100001;
rgb[6675] = 24'b001011110011011000110010;
rgb[6676] = 24'b001111110100100001000011;
rgb[6677] = 24'b010011110101101001010100;
rgb[6678] = 24'b010111110110110001100101;
rgb[6679] = 24'b011011110111111001110110;
rgb[6680] = 24'b100000001000111110000111;
rgb[6681] = 24'b100100101001111110011000;
rgb[6682] = 24'b101001001010111110101001;
rgb[6683] = 24'b101101101011111110111010;
rgb[6684] = 24'b110010001100111111001011;
rgb[6685] = 24'b110110101101111111011100;
rgb[6686] = 24'b111011001110111111101101;
rgb[6687] = 24'b111111111111111111111111;
rgb[6688] = 24'b000000000000000000000000;
rgb[6689] = 24'b000011100001001100010000;
rgb[6690] = 24'b000111010010011000100001;
rgb[6691] = 24'b001011000011100100110010;
rgb[6692] = 24'b001110100100110101000011;
rgb[6693] = 24'b010010010110000001010100;
rgb[6694] = 24'b010110000111001101100101;
rgb[6695] = 24'b011001111000011001110110;
rgb[6696] = 24'b011110001001011110000111;
rgb[6697] = 24'b100010111010011010011000;
rgb[6698] = 24'b100111101011010110101001;
rgb[6699] = 24'b101100011100010010111010;
rgb[6700] = 24'b110001011101001011001011;
rgb[6701] = 24'b110110001110000111011100;
rgb[6702] = 24'b111010111111000011101101;
rgb[6703] = 24'b111111111111111111111111;
rgb[6704] = 24'b000000000000000000000000;
rgb[6705] = 24'b000011010001010000010000;
rgb[6706] = 24'b000110110010100000100001;
rgb[6707] = 24'b001010000011110100110010;
rgb[6708] = 24'b001101100101000101000011;
rgb[6709] = 24'b010001000110010101010100;
rgb[6710] = 24'b010100010111101001100101;
rgb[6711] = 24'b010111111000111001110101;
rgb[6712] = 24'b011100001001111110000110;
rgb[6713] = 24'b100001001010110110011000;
rgb[6714] = 24'b100110001011101110101001;
rgb[6715] = 24'b101011011100100010111010;
rgb[6716] = 24'b110000011101011011001011;
rgb[6717] = 24'b110101101110001111011100;
rgb[6718] = 24'b111010101111000111101101;
rgb[6719] = 24'b111111111111111111111111;
rgb[6720] = 24'b000000000000000000000000;
rgb[6721] = 24'b000011000001010100010000;
rgb[6722] = 24'b000110000010101100100001;
rgb[6723] = 24'b001001010100000000110010;
rgb[6724] = 24'b001100010101011001000011;
rgb[6725] = 24'b001111100110101101010011;
rgb[6726] = 24'b010010101000000101100100;
rgb[6727] = 24'b010101111001011001110101;
rgb[6728] = 24'b011010001010011110000110;
rgb[6729] = 24'b011111011011010010010111;
rgb[6730] = 24'b100100111100000010101000;
rgb[6731] = 24'b101010001100110110111010;
rgb[6732] = 24'b101111101101100111001011;
rgb[6733] = 24'b110100111110011011011100;
rgb[6734] = 24'b111010011111001011101101;
rgb[6735] = 24'b111111111111111111111111;
rgb[6736] = 24'b000000000000000000000000;
rgb[6737] = 24'b000010110001011000010000;
rgb[6738] = 24'b000101100010110100100001;
rgb[6739] = 24'b001000100100010000110010;
rgb[6740] = 24'b001011010101101001000010;
rgb[6741] = 24'b001110000111000101010011;
rgb[6742] = 24'b010001001000100001100100;
rgb[6743] = 24'b010011111001111001110101;
rgb[6744] = 24'b011000001010111110000110;
rgb[6745] = 24'b011101101011101110010111;
rgb[6746] = 24'b100011011100011010101000;
rgb[6747] = 24'b101001001101000110111001;
rgb[6748] = 24'b101110111101110111001011;
rgb[6749] = 24'b110100011110100011011100;
rgb[6750] = 24'b111010001111001111101101;
rgb[6751] = 24'b111111111111111111111111;
rgb[6752] = 24'b000000000000000000000000;
rgb[6753] = 24'b000010100001011100010000;
rgb[6754] = 24'b000101000010111100100001;
rgb[6755] = 24'b000111100100011100110010;
rgb[6756] = 24'b001010000101111101000010;
rgb[6757] = 24'b001100110111011001010011;
rgb[6758] = 24'b001111011000111001100100;
rgb[6759] = 24'b010001111010011001110100;
rgb[6760] = 24'b010110001011011110000101;
rgb[6761] = 24'b011100001100000110010111;
rgb[6762] = 24'b100001111100110010101000;
rgb[6763] = 24'b100111111101011010111001;
rgb[6764] = 24'b101101111110000011001011;
rgb[6765] = 24'b110011111110101011011100;
rgb[6766] = 24'b111001111111010011101101;
rgb[6767] = 24'b111111111111111011111111;
rgb[6768] = 24'b000000000000000000000000;
rgb[6769] = 24'b000010010001100000010000;
rgb[6770] = 24'b000100100011000100100001;
rgb[6771] = 24'b000110110100101000110001;
rgb[6772] = 24'b001001000110001101000010;
rgb[6773] = 24'b001011010111110001010011;
rgb[6774] = 24'b001101101001010101100011;
rgb[6775] = 24'b001111111010111001110100;
rgb[6776] = 24'b010100001011111110000101;
rgb[6777] = 24'b011010011100100010010110;
rgb[6778] = 24'b100000101101000110101000;
rgb[6779] = 24'b100110111101101010111001;
rgb[6780] = 24'b101101001110001111001010;
rgb[6781] = 24'b110011011110110011011100;
rgb[6782] = 24'b111001101111010111101101;
rgb[6783] = 24'b111111111111111111111111;
rgb[6784] = 24'b000000000000000000000000;
rgb[6785] = 24'b000001110001101000010000;
rgb[6786] = 24'b000011110011010000100001;
rgb[6787] = 24'b000101110100111000110001;
rgb[6788] = 24'b000111110110100001000010;
rgb[6789] = 24'b001001111000001001010010;
rgb[6790] = 24'b001011111001110001100011;
rgb[6791] = 24'b001101111011011001110011;
rgb[6792] = 24'b010010001100011110000100;
rgb[6793] = 24'b011000101100111110010110;
rgb[6794] = 24'b011111001101011110100111;
rgb[6795] = 24'b100101101101111110111001;
rgb[6796] = 24'b101100001110011111001010;
rgb[6797] = 24'b110010101110111111011100;
rgb[6798] = 24'b111001001111011111101101;
rgb[6799] = 24'b111111111111111011111111;
rgb[6800] = 24'b000000000000000000000000;
rgb[6801] = 24'b000001100001101100010000;
rgb[6802] = 24'b000011010011011000100001;
rgb[6803] = 24'b000101000101000100110001;
rgb[6804] = 24'b000110110110110001000010;
rgb[6805] = 24'b001000011000100001010010;
rgb[6806] = 24'b001010001010001101100011;
rgb[6807] = 24'b001011111011111001110011;
rgb[6808] = 24'b010000001100111110000100;
rgb[6809] = 24'b010110111101011010010110;
rgb[6810] = 24'b011101101101110110100111;
rgb[6811] = 24'b100100101110001110111001;
rgb[6812] = 24'b101011011110101011001010;
rgb[6813] = 24'b110010001111000111011100;
rgb[6814] = 24'b111000111111100011101101;
rgb[6815] = 24'b111111111111111111111111;
rgb[6816] = 24'b000000000000000000000000;
rgb[6817] = 24'b000001010001110000010000;
rgb[6818] = 24'b000010110011100000100000;
rgb[6819] = 24'b000100010101010100110001;
rgb[6820] = 24'b000101100111000101000001;
rgb[6821] = 24'b000111001000110101010010;
rgb[6822] = 24'b001000101010101001100010;
rgb[6823] = 24'b001001111100011001110011;
rgb[6824] = 24'b001110001101011110000100;
rgb[6825] = 24'b010101001101110110010101;
rgb[6826] = 24'b011100011110001010100111;
rgb[6827] = 24'b100011011110100010111000;
rgb[6828] = 24'b101010101110111011001010;
rgb[6829] = 24'b110001101111001111011011;
rgb[6830] = 24'b111000101111100111101101;
rgb[6831] = 24'b111111111111111011111111;
rgb[6832] = 24'b000000000000000000000000;
rgb[6833] = 24'b000001000001110100010000;
rgb[6834] = 24'b000010010011101000100000;
rgb[6835] = 24'b000011010101100000110001;
rgb[6836] = 24'b000100100111010101000001;
rgb[6837] = 24'b000101101001001101010010;
rgb[6838] = 24'b000110111011000001100010;
rgb[6839] = 24'b000111111100111001110010;
rgb[6840] = 24'b001100001101111110000011;
rgb[6841] = 24'b010011101110001110010101;
rgb[6842] = 24'b011010111110100010100111;
rgb[6843] = 24'b100010011110110010111000;
rgb[6844] = 24'b101001101111000111001010;
rgb[6845] = 24'b110001001111010111011011;
rgb[6846] = 24'b111000011111101011101101;
rgb[6847] = 24'b111111111111111111111111;
rgb[6848] = 24'b000000000000000000000000;
rgb[6849] = 24'b000000110001111000010000;
rgb[6850] = 24'b000001100011110100100000;
rgb[6851] = 24'b000010100101101100110001;
rgb[6852] = 24'b000011010111101001000001;
rgb[6853] = 24'b000100001001100101010001;
rgb[6854] = 24'b000101001011011101100010;
rgb[6855] = 24'b000101111101011001110010;
rgb[6856] = 24'b001010001110011110000011;
rgb[6857] = 24'b010001111110101010010101;
rgb[6858] = 24'b011001011110111010100110;
rgb[6859] = 24'b100001001111000110111000;
rgb[6860] = 24'b101000111111010011001010;
rgb[6861] = 24'b110000011111100011011011;
rgb[6862] = 24'b111000001111101111101101;
rgb[6863] = 24'b111111111111111111111111;
rgb[6864] = 24'b000000000000000000000000;
rgb[6865] = 24'b000000100001111100010000;
rgb[6866] = 24'b000001000011111100100000;
rgb[6867] = 24'b000001100101111100110000;
rgb[6868] = 24'b000010010111111001000001;
rgb[6869] = 24'b000010111001111001010001;
rgb[6870] = 24'b000011011011111001100001;
rgb[6871] = 24'b000011111101111001110010;
rgb[6872] = 24'b001000001110111110000011;
rgb[6873] = 24'b010000001111000110010100;
rgb[6874] = 24'b011000001111001110100110;
rgb[6875] = 24'b100000001111010110111000;
rgb[6876] = 24'b100111111111100011001001;
rgb[6877] = 24'b101111111111101011011011;
rgb[6878] = 24'b110111111111110011101101;
rgb[6879] = 24'b111111111111111111111111;
rgb[6880] = 24'b000000000000000000000000;
rgb[6881] = 24'b000000010010000000010000;
rgb[6882] = 24'b000000100100000100100000;
rgb[6883] = 24'b000000110110001000110000;
rgb[6884] = 24'b000001001000001101000000;
rgb[6885] = 24'b000001011010010001010001;
rgb[6886] = 24'b000001101100010101100001;
rgb[6887] = 24'b000001111110011001110001;
rgb[6888] = 24'b000110001111011110000010;
rgb[6889] = 24'b001110011111100010010100;
rgb[6890] = 24'b010110101111100110100110;
rgb[6891] = 24'b011110111111101010110111;
rgb[6892] = 24'b100111001111101111001001;
rgb[6893] = 24'b101111011111110011011011;
rgb[6894] = 24'b110111101111110111101101;
rgb[6895] = 24'b111111111111111111111111;
rgb[6896] = 24'b000000000000000000000000;
rgb[6897] = 24'b000000000010001000010000;
rgb[6898] = 24'b000000000100010000100000;
rgb[6899] = 24'b000000000110011000110000;
rgb[6900] = 24'b000000001000100001000000;
rgb[6901] = 24'b000000001010101001010000;
rgb[6902] = 24'b000000001100110001100001;
rgb[6903] = 24'b000000001110111001110001;
rgb[6904] = 24'b000100011111111010000010;
rgb[6905] = 24'b001100101111111110010100;
rgb[6906] = 24'b010101011111111010100101;
rgb[6907] = 24'b011101101111111110110111;
rgb[6908] = 24'b100110011111111111001001;
rgb[6909] = 24'b101110111111111111011011;
rgb[6910] = 24'b110111011111111111101101;
rgb[6911] = 24'b111111111111111111111111;
rgb[6912] = 24'b000000000000000000000000;
rgb[6913] = 24'b000100010001000100010001;
rgb[6914] = 24'b001000100010001000100010;
rgb[6915] = 24'b001100110011001100110011;
rgb[6916] = 24'b010001000100010001000100;
rgb[6917] = 24'b010101010101010101010101;
rgb[6918] = 24'b011001100110011001100110;
rgb[6919] = 24'b011101110111011101110111;
rgb[6920] = 24'b100010001000100010001000;
rgb[6921] = 24'b100110011001100110011001;
rgb[6922] = 24'b101010101010101010101010;
rgb[6923] = 24'b101110111011101110111011;
rgb[6924] = 24'b110011001100110011001100;
rgb[6925] = 24'b110111011101110111011101;
rgb[6926] = 24'b111011101110111011101110;
rgb[6927] = 24'b111111111111111111111111;
rgb[6928] = 24'b000000000000000000000000;
rgb[6929] = 24'b000011110001001000010001;
rgb[6930] = 24'b000111110010010000100010;
rgb[6931] = 24'b001011110011011000110011;
rgb[6932] = 24'b001111110100100001000100;
rgb[6933] = 24'b010011110101101001010101;
rgb[6934] = 24'b010111110110110001100110;
rgb[6935] = 24'b011011110111111001111000;
rgb[6936] = 24'b100000001000111110001001;
rgb[6937] = 24'b100100101001111110011001;
rgb[6938] = 24'b101001001010111110101010;
rgb[6939] = 24'b101101101011111110111011;
rgb[6940] = 24'b110010001100111111001100;
rgb[6941] = 24'b110110101101111111011101;
rgb[6942] = 24'b111011001110111111101110;
rgb[6943] = 24'b111111111111111111111111;
rgb[6944] = 24'b000000000000000000000000;
rgb[6945] = 24'b000011100001001100010001;
rgb[6946] = 24'b000111010010011000100010;
rgb[6947] = 24'b001011000011100100110011;
rgb[6948] = 24'b001110100100110101000101;
rgb[6949] = 24'b010010010110000001010110;
rgb[6950] = 24'b010110000111001101100111;
rgb[6951] = 24'b011001111000011001111001;
rgb[6952] = 24'b011110001001011110001010;
rgb[6953] = 24'b100010111010011010011010;
rgb[6954] = 24'b100111101011010110101011;
rgb[6955] = 24'b101100011100010010111100;
rgb[6956] = 24'b110001011101001011001100;
rgb[6957] = 24'b110110001110000111011101;
rgb[6958] = 24'b111010111111000011101110;
rgb[6959] = 24'b111111111111111111111111;
rgb[6960] = 24'b000000000000000000000000;
rgb[6961] = 24'b000011010001010000010001;
rgb[6962] = 24'b000110110010100000100010;
rgb[6963] = 24'b001010000011110100110100;
rgb[6964] = 24'b001101100101000101000101;
rgb[6965] = 24'b010001000110010101010111;
rgb[6966] = 24'b010100010111101001101000;
rgb[6967] = 24'b010111111000111001111010;
rgb[6968] = 24'b011100001001111110001011;
rgb[6969] = 24'b100001001010110110011011;
rgb[6970] = 24'b100110001011101110101100;
rgb[6971] = 24'b101011011100100010111100;
rgb[6972] = 24'b110000011101011011001101;
rgb[6973] = 24'b110101101110001111011101;
rgb[6974] = 24'b111010101111000111101110;
rgb[6975] = 24'b111111111111111111111111;
rgb[6976] = 24'b000000000000000000000000;
rgb[6977] = 24'b000011000001010100010001;
rgb[6978] = 24'b000110000010101100100011;
rgb[6979] = 24'b001001010100000000110100;
rgb[6980] = 24'b001100010101011001000110;
rgb[6981] = 24'b001111100110101101011000;
rgb[6982] = 24'b010010101000000101101001;
rgb[6983] = 24'b010101111001011001111011;
rgb[6984] = 24'b011010001010011110001100;
rgb[6985] = 24'b011111011011010010011100;
rgb[6986] = 24'b100100111100000010101101;
rgb[6987] = 24'b101010001100110110111101;
rgb[6988] = 24'b101111101101100111001101;
rgb[6989] = 24'b110100111110011011011110;
rgb[6990] = 24'b111010011111001011101110;
rgb[6991] = 24'b111111111111111111111111;
rgb[6992] = 24'b000000000000000000000000;
rgb[6993] = 24'b000010110001011000010001;
rgb[6994] = 24'b000101100010110100100011;
rgb[6995] = 24'b001000100100010000110101;
rgb[6996] = 24'b001011010101101001000111;
rgb[6997] = 24'b001110000111000101011001;
rgb[6998] = 24'b010001001000100001101010;
rgb[6999] = 24'b010011111001111001111100;
rgb[7000] = 24'b011000001010111110001101;
rgb[7001] = 24'b011101101011101110011101;
rgb[7002] = 24'b100011011100011010101110;
rgb[7003] = 24'b101001001101000110111110;
rgb[7004] = 24'b101110111101110111001110;
rgb[7005] = 24'b110100011110100011011110;
rgb[7006] = 24'b111010001111001111101110;
rgb[7007] = 24'b111111111111111111111111;
rgb[7008] = 24'b000000000000000000000000;
rgb[7009] = 24'b000010100001011100010001;
rgb[7010] = 24'b000101000010111100100011;
rgb[7011] = 24'b000111100100011100110101;
rgb[7012] = 24'b001010000101111101000111;
rgb[7013] = 24'b001100110111011001011001;
rgb[7014] = 24'b001111011000111001101011;
rgb[7015] = 24'b010001111010011001111101;
rgb[7016] = 24'b010110001011011110001110;
rgb[7017] = 24'b011100001100000110011110;
rgb[7018] = 24'b100001111100110010101110;
rgb[7019] = 24'b100111111101011010111110;
rgb[7020] = 24'b101101111110000011001110;
rgb[7021] = 24'b110011111110101011011110;
rgb[7022] = 24'b111001111111010011101110;
rgb[7023] = 24'b111111111111111011111110;
rgb[7024] = 24'b000000000000000000000000;
rgb[7025] = 24'b000010010001100000010010;
rgb[7026] = 24'b000100100011000100100100;
rgb[7027] = 24'b000110110100101000110110;
rgb[7028] = 24'b001001000110001101001000;
rgb[7029] = 24'b001011010111110001011010;
rgb[7030] = 24'b001101101001010101101100;
rgb[7031] = 24'b001111111010111001111110;
rgb[7032] = 24'b010100001011111110001111;
rgb[7033] = 24'b011010011100100010011111;
rgb[7034] = 24'b100000101101000110101111;
rgb[7035] = 24'b100110111101101010111111;
rgb[7036] = 24'b101101001110001111001111;
rgb[7037] = 24'b110011011110110011011111;
rgb[7038] = 24'b111001101111010111101111;
rgb[7039] = 24'b111111111111111111111111;
rgb[7040] = 24'b000000000000000000000000;
rgb[7041] = 24'b000001110001101000010010;
rgb[7042] = 24'b000011110011010000100100;
rgb[7043] = 24'b000101110100111000110110;
rgb[7044] = 24'b000111110110100001001001;
rgb[7045] = 24'b001001111000001001011011;
rgb[7046] = 24'b001011111001110001101101;
rgb[7047] = 24'b001101111011011010000000;
rgb[7048] = 24'b010010001100011110010001;
rgb[7049] = 24'b011000101100111110100000;
rgb[7050] = 24'b011111001101011110110000;
rgb[7051] = 24'b100101101101111111000000;
rgb[7052] = 24'b101100001110011111001111;
rgb[7053] = 24'b110010101110111111011111;
rgb[7054] = 24'b111001001111011111101111;
rgb[7055] = 24'b111111111111111011111110;
rgb[7056] = 24'b000000000000000000000000;
rgb[7057] = 24'b000001100001101100010010;
rgb[7058] = 24'b000011010011011000100100;
rgb[7059] = 24'b000101000101000100110111;
rgb[7060] = 24'b000110110110110001001001;
rgb[7061] = 24'b001000011000100001011100;
rgb[7062] = 24'b001010001010001101101110;
rgb[7063] = 24'b001011111011111010000001;
rgb[7064] = 24'b010000001100111110010010;
rgb[7065] = 24'b010110111101011010100001;
rgb[7066] = 24'b011101101101110110110001;
rgb[7067] = 24'b100100101110001111000000;
rgb[7068] = 24'b101011011110101011010000;
rgb[7069] = 24'b110010001111000111011111;
rgb[7070] = 24'b111000111111100011101111;
rgb[7071] = 24'b111111111111111111111111;
rgb[7072] = 24'b000000000000000000000000;
rgb[7073] = 24'b000001010001110000010010;
rgb[7074] = 24'b000010110011100000100101;
rgb[7075] = 24'b000100010101010100110111;
rgb[7076] = 24'b000101100111000101001010;
rgb[7077] = 24'b000111001000110101011101;
rgb[7078] = 24'b001000101010101001101111;
rgb[7079] = 24'b001001111100011010000010;
rgb[7080] = 24'b001110001101011110010011;
rgb[7081] = 24'b010101001101110110100010;
rgb[7082] = 24'b011100011110001010110010;
rgb[7083] = 24'b100011011110100011000001;
rgb[7084] = 24'b101010101110111011010000;
rgb[7085] = 24'b110001101111001111100000;
rgb[7086] = 24'b111000101111100111101111;
rgb[7087] = 24'b111111111111111011111110;
rgb[7088] = 24'b000000000000000000000000;
rgb[7089] = 24'b000001000001110100010010;
rgb[7090] = 24'b000010010011101000100101;
rgb[7091] = 24'b000011010101100000111000;
rgb[7092] = 24'b000100100111010101001011;
rgb[7093] = 24'b000101101001001101011101;
rgb[7094] = 24'b000110111011000001110000;
rgb[7095] = 24'b000111111100111010000011;
rgb[7096] = 24'b001100001101111110010100;
rgb[7097] = 24'b010011101110001110100011;
rgb[7098] = 24'b011010111110100010110010;
rgb[7099] = 24'b100010011110110011000010;
rgb[7100] = 24'b101001101111000111010001;
rgb[7101] = 24'b110001001111010111100000;
rgb[7102] = 24'b111000011111101011101111;
rgb[7103] = 24'b111111111111111111111111;
rgb[7104] = 24'b000000000000000000000000;
rgb[7105] = 24'b000000110001111000010010;
rgb[7106] = 24'b000001100011110100100101;
rgb[7107] = 24'b000010100101101100111000;
rgb[7108] = 24'b000011010111101001001011;
rgb[7109] = 24'b000100001001100101011110;
rgb[7110] = 24'b000101001011011101110001;
rgb[7111] = 24'b000101111101011010000100;
rgb[7112] = 24'b001010001110011110010101;
rgb[7113] = 24'b010001111110101010100100;
rgb[7114] = 24'b011001011110111010110011;
rgb[7115] = 24'b100001001111000111000010;
rgb[7116] = 24'b101000111111010011010001;
rgb[7117] = 24'b110000011111100011100000;
rgb[7118] = 24'b111000001111101111101111;
rgb[7119] = 24'b111111111111111111111111;
rgb[7120] = 24'b000000000000000000000000;
rgb[7121] = 24'b000000100001111100010011;
rgb[7122] = 24'b000001000011111100100110;
rgb[7123] = 24'b000001100101111100111001;
rgb[7124] = 24'b000010010111111001001100;
rgb[7125] = 24'b000010111001111001011111;
rgb[7126] = 24'b000011011011111001110010;
rgb[7127] = 24'b000011111101111010000101;
rgb[7128] = 24'b001000001110111110010110;
rgb[7129] = 24'b010000001111000110100101;
rgb[7130] = 24'b011000001111001110110100;
rgb[7131] = 24'b100000001111010111000011;
rgb[7132] = 24'b100111111111100011010010;
rgb[7133] = 24'b101111111111101011100001;
rgb[7134] = 24'b110111111111110011110000;
rgb[7135] = 24'b111111111111111111111111;
rgb[7136] = 24'b000000000000000000000000;
rgb[7137] = 24'b000000010010000000010011;
rgb[7138] = 24'b000000100100000100100110;
rgb[7139] = 24'b000000110110001000111001;
rgb[7140] = 24'b000001001000001101001101;
rgb[7141] = 24'b000001011010010001100000;
rgb[7142] = 24'b000001101100010101110011;
rgb[7143] = 24'b000001111110011010000110;
rgb[7144] = 24'b000110001111011110010111;
rgb[7145] = 24'b001110011111100010100110;
rgb[7146] = 24'b010110101111100110110101;
rgb[7147] = 24'b011110111111101011000100;
rgb[7148] = 24'b100111001111101111010010;
rgb[7149] = 24'b101111011111110011100001;
rgb[7150] = 24'b110111101111110111110000;
rgb[7151] = 24'b111111111111111111111111;
rgb[7152] = 24'b000000000000000000000000;
rgb[7153] = 24'b000000000010001000010011;
rgb[7154] = 24'b000000000100010000100110;
rgb[7155] = 24'b000000000110011000111010;
rgb[7156] = 24'b000000001000100001001101;
rgb[7157] = 24'b000000001010101001100001;
rgb[7158] = 24'b000000001100110001110100;
rgb[7159] = 24'b000000001110111010001000;
rgb[7160] = 24'b000100011111111010011001;
rgb[7161] = 24'b001100101111111110100111;
rgb[7162] = 24'b010101011111111010110110;
rgb[7163] = 24'b011101101111111111000100;
rgb[7164] = 24'b100110011111111111010011;
rgb[7165] = 24'b101110111111111111100001;
rgb[7166] = 24'b110111011111111111110000;
rgb[7167] = 24'b111111111111111111111111;
rgb[7168] = 24'b000000000000000000000000;
rgb[7169] = 24'b000100010001000100010001;
rgb[7170] = 24'b001000100010001000100010;
rgb[7171] = 24'b001100110011001100110011;
rgb[7172] = 24'b010001000100010001000100;
rgb[7173] = 24'b010101010101010101010101;
rgb[7174] = 24'b011001100110011001100110;
rgb[7175] = 24'b011101110111011101110111;
rgb[7176] = 24'b100010001000100010001000;
rgb[7177] = 24'b100110011001100110011001;
rgb[7178] = 24'b101010101010101010101010;
rgb[7179] = 24'b101110111011101110111011;
rgb[7180] = 24'b110011001100110011001100;
rgb[7181] = 24'b110111011101110111011101;
rgb[7182] = 24'b111011101110111011101110;
rgb[7183] = 24'b111111111111111111111111;
rgb[7184] = 24'b000000000000000000000000;
rgb[7185] = 24'b000011110001001000010001;
rgb[7186] = 24'b000111110010010000100010;
rgb[7187] = 24'b001011110011011000110100;
rgb[7188] = 24'b001111110100100001000101;
rgb[7189] = 24'b010011110101101001010110;
rgb[7190] = 24'b010111110110110001101000;
rgb[7191] = 24'b011011110111111001111001;
rgb[7192] = 24'b100000001000111110001010;
rgb[7193] = 24'b100100101001111110011011;
rgb[7194] = 24'b101001001010111110101011;
rgb[7195] = 24'b101101101011111110111100;
rgb[7196] = 24'b110010001100111111001101;
rgb[7197] = 24'b110110101101111111011101;
rgb[7198] = 24'b111011001110111111101110;
rgb[7199] = 24'b111111111111111111111111;
rgb[7200] = 24'b000000000000000000000000;
rgb[7201] = 24'b000011100001001100010001;
rgb[7202] = 24'b000111010010011000100011;
rgb[7203] = 24'b001011000011100100110101;
rgb[7204] = 24'b001110100100110101000111;
rgb[7205] = 24'b010010010110000001011000;
rgb[7206] = 24'b010110000111001101101010;
rgb[7207] = 24'b011001111000011001111100;
rgb[7208] = 24'b011110001001011110001101;
rgb[7209] = 24'b100010111010011010011101;
rgb[7210] = 24'b100111101011010110101101;
rgb[7211] = 24'b101100011100010010111110;
rgb[7212] = 24'b110001011101001011001110;
rgb[7213] = 24'b110110001110000111011110;
rgb[7214] = 24'b111010111111000011101110;
rgb[7215] = 24'b111111111111111111111111;
rgb[7216] = 24'b000000000000000000000000;
rgb[7217] = 24'b000011010001010000010010;
rgb[7218] = 24'b000110110010100000100100;
rgb[7219] = 24'b001010000011110100110110;
rgb[7220] = 24'b001101100101000101001000;
rgb[7221] = 24'b010001000110010101011010;
rgb[7222] = 24'b010100010111101001101100;
rgb[7223] = 24'b010111111000111001111110;
rgb[7224] = 24'b011100001001111110001111;
rgb[7225] = 24'b100001001010110110011111;
rgb[7226] = 24'b100110001011101110101111;
rgb[7227] = 24'b101011011100100010111111;
rgb[7228] = 24'b110000011101011011001111;
rgb[7229] = 24'b110101101110001111011111;
rgb[7230] = 24'b111010101111000111101111;
rgb[7231] = 24'b111111111111111111111111;
rgb[7232] = 24'b000000000000000000000000;
rgb[7233] = 24'b000011000001010100010010;
rgb[7234] = 24'b000110000010101100100101;
rgb[7235] = 24'b001001010100000000110111;
rgb[7236] = 24'b001100010101011001001010;
rgb[7237] = 24'b001111100110101101011100;
rgb[7238] = 24'b010010101000000101101111;
rgb[7239] = 24'b010101111001011010000001;
rgb[7240] = 24'b011010001010011110010010;
rgb[7241] = 24'b011111011011010010100010;
rgb[7242] = 24'b100100111100000010110001;
rgb[7243] = 24'b101010001100110111000001;
rgb[7244] = 24'b101111101101100111010000;
rgb[7245] = 24'b110100111110011011100000;
rgb[7246] = 24'b111010011111001011101111;
rgb[7247] = 24'b111111111111111111111111;
rgb[7248] = 24'b000000000000000000000000;
rgb[7249] = 24'b000010110001011000010010;
rgb[7250] = 24'b000101100010110100100101;
rgb[7251] = 24'b001000100100010000111000;
rgb[7252] = 24'b001011010101101001001011;
rgb[7253] = 24'b001110000111000101011110;
rgb[7254] = 24'b010001001000100001110001;
rgb[7255] = 24'b010011111001111010000100;
rgb[7256] = 24'b011000001010111110010101;
rgb[7257] = 24'b011101101011101110100100;
rgb[7258] = 24'b100011011100011010110011;
rgb[7259] = 24'b101001001101000111000010;
rgb[7260] = 24'b101110111101110111010001;
rgb[7261] = 24'b110100011110100011100000;
rgb[7262] = 24'b111010001111001111101111;
rgb[7263] = 24'b111111111111111111111111;
rgb[7264] = 24'b000000000000000000000000;
rgb[7265] = 24'b000010100001011100010011;
rgb[7266] = 24'b000101000010111100100110;
rgb[7267] = 24'b000111100100011100111001;
rgb[7268] = 24'b001010000101111101001101;
rgb[7269] = 24'b001100110111011001100000;
rgb[7270] = 24'b001111011000111001110011;
rgb[7271] = 24'b010001111010011010000110;
rgb[7272] = 24'b010110001011011110010111;
rgb[7273] = 24'b011100001100000110100110;
rgb[7274] = 24'b100001111100110010110101;
rgb[7275] = 24'b100111111101011011000100;
rgb[7276] = 24'b101101111110000011010010;
rgb[7277] = 24'b110011111110101011100001;
rgb[7278] = 24'b111001111111010011110000;
rgb[7279] = 24'b111111111111111011111110;
rgb[7280] = 24'b000000000000000000000000;
rgb[7281] = 24'b000010010001100000010011;
rgb[7282] = 24'b000100100011000100100111;
rgb[7283] = 24'b000110110100101000111010;
rgb[7284] = 24'b001001000110001101001110;
rgb[7285] = 24'b001011010111110001100010;
rgb[7286] = 24'b001101101001010101110101;
rgb[7287] = 24'b001111111010111010001001;
rgb[7288] = 24'b010100001011111110011010;
rgb[7289] = 24'b011010011100100010101000;
rgb[7290] = 24'b100000101101000110110111;
rgb[7291] = 24'b100110111101101011000101;
rgb[7292] = 24'b101101001110001111010011;
rgb[7293] = 24'b110011011110110011100010;
rgb[7294] = 24'b111001101111010111110000;
rgb[7295] = 24'b111111111111111111111111;
rgb[7296] = 24'b000000000000000000000000;
rgb[7297] = 24'b000001110001101000010100;
rgb[7298] = 24'b000011110011010000101000;
rgb[7299] = 24'b000101110100111000111100;
rgb[7300] = 24'b000111110110100001010000;
rgb[7301] = 24'b001001111000001001100100;
rgb[7302] = 24'b001011111001110001111000;
rgb[7303] = 24'b001101111011011010001100;
rgb[7304] = 24'b010010001100011110011101;
rgb[7305] = 24'b011000101100111110101011;
rgb[7306] = 24'b011111001101011110111001;
rgb[7307] = 24'b100101101101111111000111;
rgb[7308] = 24'b101100001110011111010101;
rgb[7309] = 24'b110010101110111111100011;
rgb[7310] = 24'b111001001111011111110001;
rgb[7311] = 24'b111111111111111011111110;
rgb[7312] = 24'b000000000000000000000000;
rgb[7313] = 24'b000001100001101100010100;
rgb[7314] = 24'b000011010011011000101000;
rgb[7315] = 24'b000101000101000100111101;
rgb[7316] = 24'b000110110110110001010001;
rgb[7317] = 24'b001000011000100001100101;
rgb[7318] = 24'b001010001010001101111010;
rgb[7319] = 24'b001011111011111010001110;
rgb[7320] = 24'b010000001100111110011111;
rgb[7321] = 24'b010110111101011010101101;
rgb[7322] = 24'b011101101101110110111011;
rgb[7323] = 24'b100100101110001111001000;
rgb[7324] = 24'b101011011110101011010110;
rgb[7325] = 24'b110010001111000111100011;
rgb[7326] = 24'b111000111111100011110001;
rgb[7327] = 24'b111111111111111111111111;
rgb[7328] = 24'b000000000000000000000000;
rgb[7329] = 24'b000001010001110000010100;
rgb[7330] = 24'b000010110011100000101001;
rgb[7331] = 24'b000100010101010100111110;
rgb[7332] = 24'b000101100111000101010011;
rgb[7333] = 24'b000111001000110101100111;
rgb[7334] = 24'b001000101010101001111100;
rgb[7335] = 24'b001001111100011010010001;
rgb[7336] = 24'b001110001101011110100010;
rgb[7337] = 24'b010101001101110110101111;
rgb[7338] = 24'b011100011110001010111100;
rgb[7339] = 24'b100011011110100011001010;
rgb[7340] = 24'b101010101110111011010111;
rgb[7341] = 24'b110001101111001111100100;
rgb[7342] = 24'b111000101111100111110001;
rgb[7343] = 24'b111111111111111011111110;
rgb[7344] = 24'b000000000000000000000000;
rgb[7345] = 24'b000001000001110100010101;
rgb[7346] = 24'b000010010011101000101010;
rgb[7347] = 24'b000011010101100000111111;
rgb[7348] = 24'b000100100111010101010100;
rgb[7349] = 24'b000101101001001101101001;
rgb[7350] = 24'b000110111011000001111110;
rgb[7351] = 24'b000111111100111010010100;
rgb[7352] = 24'b001100001101111110100101;
rgb[7353] = 24'b010011101110001110110001;
rgb[7354] = 24'b011010111110100010111110;
rgb[7355] = 24'b100010011110110011001011;
rgb[7356] = 24'b101001101111000111011000;
rgb[7357] = 24'b110001001111010111100101;
rgb[7358] = 24'b111000011111101011110010;
rgb[7359] = 24'b111111111111111111111111;
rgb[7360] = 24'b000000000000000000000000;
rgb[7361] = 24'b000000110001111000010101;
rgb[7362] = 24'b000001100011110100101011;
rgb[7363] = 24'b000010100101101101000000;
rgb[7364] = 24'b000011010111101001010110;
rgb[7365] = 24'b000100001001100101101011;
rgb[7366] = 24'b000101001011011110000001;
rgb[7367] = 24'b000101111101011010010110;
rgb[7368] = 24'b001010001110011110100111;
rgb[7369] = 24'b010001111110101010110100;
rgb[7370] = 24'b011001011110111011000000;
rgb[7371] = 24'b100001001111000111001101;
rgb[7372] = 24'b101000111111010011011001;
rgb[7373] = 24'b110000011111100011100110;
rgb[7374] = 24'b111000001111101111110010;
rgb[7375] = 24'b111111111111111111111111;
rgb[7376] = 24'b000000000000000000000000;
rgb[7377] = 24'b000000100001111100010101;
rgb[7378] = 24'b000001000011111100101011;
rgb[7379] = 24'b000001100101111101000001;
rgb[7380] = 24'b000010010111111001010111;
rgb[7381] = 24'b000010111001111001101101;
rgb[7382] = 24'b000011011011111010000011;
rgb[7383] = 24'b000011111101111010011001;
rgb[7384] = 24'b001000001110111110101010;
rgb[7385] = 24'b010000001111000110110110;
rgb[7386] = 24'b011000001111001111000010;
rgb[7387] = 24'b100000001111010111001110;
rgb[7388] = 24'b100111111111100011011010;
rgb[7389] = 24'b101111111111101011100110;
rgb[7390] = 24'b110111111111110011110010;
rgb[7391] = 24'b111111111111111111111111;
rgb[7392] = 24'b000000000000000000000000;
rgb[7393] = 24'b000000010010000000010110;
rgb[7394] = 24'b000000100100000100101100;
rgb[7395] = 24'b000000110110001001000010;
rgb[7396] = 24'b000001001000001101011001;
rgb[7397] = 24'b000001011010010001101111;
rgb[7398] = 24'b000001101100010110000101;
rgb[7399] = 24'b000001111110011010011100;
rgb[7400] = 24'b000110001111011110101101;
rgb[7401] = 24'b001110011111100010111000;
rgb[7402] = 24'b010110101111100111000100;
rgb[7403] = 24'b011110111111101011010000;
rgb[7404] = 24'b100111001111101111011011;
rgb[7405] = 24'b101111011111110011100111;
rgb[7406] = 24'b110111101111110111110011;
rgb[7407] = 24'b111111111111111111111111;
rgb[7408] = 24'b000000000000000000000000;
rgb[7409] = 24'b000000000010001000010110;
rgb[7410] = 24'b000000000100010000101101;
rgb[7411] = 24'b000000000110011001000100;
rgb[7412] = 24'b000000001000100001011010;
rgb[7413] = 24'b000000001010101001110001;
rgb[7414] = 24'b000000001100110010001000;
rgb[7415] = 24'b000000001110111010011110;
rgb[7416] = 24'b000100011111111010101111;
rgb[7417] = 24'b001100101111111110111011;
rgb[7418] = 24'b010101011111111011000110;
rgb[7419] = 24'b011101101111111111010001;
rgb[7420] = 24'b100110011111111111011101;
rgb[7421] = 24'b101110111111111111101000;
rgb[7422] = 24'b110111011111111111110011;
rgb[7423] = 24'b111111111111111111111111;
rgb[7424] = 24'b000000000000000000000000;
rgb[7425] = 24'b000100010001000100010001;
rgb[7426] = 24'b001000100010001000100010;
rgb[7427] = 24'b001100110011001100110011;
rgb[7428] = 24'b010001000100010001000100;
rgb[7429] = 24'b010101010101010101010101;
rgb[7430] = 24'b011001100110011001100110;
rgb[7431] = 24'b011101110111011101110111;
rgb[7432] = 24'b100010001000100010001000;
rgb[7433] = 24'b100110011001100110011001;
rgb[7434] = 24'b101010101010101010101010;
rgb[7435] = 24'b101110111011101110111011;
rgb[7436] = 24'b110011001100110011001100;
rgb[7437] = 24'b110111011101110111011101;
rgb[7438] = 24'b111011101110111011101110;
rgb[7439] = 24'b111111111111111111111111;
rgb[7440] = 24'b000000000000000000000000;
rgb[7441] = 24'b000011110001001000010001;
rgb[7442] = 24'b000111110010010000100011;
rgb[7443] = 24'b001011110011011000110100;
rgb[7444] = 24'b001111110100100001000110;
rgb[7445] = 24'b010011110101101001010111;
rgb[7446] = 24'b010111110110110001101001;
rgb[7447] = 24'b011011110111111001111011;
rgb[7448] = 24'b100000001000111110001100;
rgb[7449] = 24'b100100101001111110011100;
rgb[7450] = 24'b101001001010111110101100;
rgb[7451] = 24'b101101101011111110111101;
rgb[7452] = 24'b110010001100111111001101;
rgb[7453] = 24'b110110101101111111011110;
rgb[7454] = 24'b111011001110111111101110;
rgb[7455] = 24'b111111111111111111111111;
rgb[7456] = 24'b000000000000000000000000;
rgb[7457] = 24'b000011100001001100010010;
rgb[7458] = 24'b000111010010011000100100;
rgb[7459] = 24'b001011000011100100110110;
rgb[7460] = 24'b001110100100110101001000;
rgb[7461] = 24'b010010010110000001011010;
rgb[7462] = 24'b010110000111001101101101;
rgb[7463] = 24'b011001111000011001111111;
rgb[7464] = 24'b011110001001011110010000;
rgb[7465] = 24'b100010111010011010100000;
rgb[7466] = 24'b100111101011010110101111;
rgb[7467] = 24'b101100011100010010111111;
rgb[7468] = 24'b110001011101001011001111;
rgb[7469] = 24'b110110001110000111011111;
rgb[7470] = 24'b111010111111000011101111;
rgb[7471] = 24'b111111111111111111111111;
rgb[7472] = 24'b000000000000000000000000;
rgb[7473] = 24'b000011010001010000010010;
rgb[7474] = 24'b000110110010100000100101;
rgb[7475] = 24'b001010000011110100111000;
rgb[7476] = 24'b001101100101000101001011;
rgb[7477] = 24'b010001000110010101011101;
rgb[7478] = 24'b010100010111101001110000;
rgb[7479] = 24'b010111111000111010000011;
rgb[7480] = 24'b011100001001111110010100;
rgb[7481] = 24'b100001001010110110100011;
rgb[7482] = 24'b100110001011101110110010;
rgb[7483] = 24'b101011011100100011000010;
rgb[7484] = 24'b110000011101011011010001;
rgb[7485] = 24'b110101101110001111100000;
rgb[7486] = 24'b111010101111000111101111;
rgb[7487] = 24'b111111111111111111111111;
rgb[7488] = 24'b000000000000000000000000;
rgb[7489] = 24'b000011000001010100010011;
rgb[7490] = 24'b000110000010101100100110;
rgb[7491] = 24'b001001010100000000111010;
rgb[7492] = 24'b001100010101011001001101;
rgb[7493] = 24'b001111100110101101100000;
rgb[7494] = 24'b010010101000000101110100;
rgb[7495] = 24'b010101111001011010000111;
rgb[7496] = 24'b011010001010011110011000;
rgb[7497] = 24'b011111011011010010100111;
rgb[7498] = 24'b100100111100000010110101;
rgb[7499] = 24'b101010001100110111000100;
rgb[7500] = 24'b101111101101100111010011;
rgb[7501] = 24'b110100111110011011100001;
rgb[7502] = 24'b111010011111001011110000;
rgb[7503] = 24'b111111111111111111111111;
rgb[7504] = 24'b000000000000000000000000;
rgb[7505] = 24'b000010110001011000010011;
rgb[7506] = 24'b000101100010110100100111;
rgb[7507] = 24'b001000100100010000111011;
rgb[7508] = 24'b001011010101101001001111;
rgb[7509] = 24'b001110000111000101100011;
rgb[7510] = 24'b010001001000100001110111;
rgb[7511] = 24'b010011111001111010001011;
rgb[7512] = 24'b011000001010111110011100;
rgb[7513] = 24'b011101101011101110101010;
rgb[7514] = 24'b100011011100011010111000;
rgb[7515] = 24'b101001001101000111000110;
rgb[7516] = 24'b101110111101110111010100;
rgb[7517] = 24'b110100011110100011100010;
rgb[7518] = 24'b111010001111001111110000;
rgb[7519] = 24'b111111111111111111111111;
rgb[7520] = 24'b000000000000000000000000;
rgb[7521] = 24'b000010100001011100010100;
rgb[7522] = 24'b000101000010111100101001;
rgb[7523] = 24'b000111100100011100111101;
rgb[7524] = 24'b001010000101111101010010;
rgb[7525] = 24'b001100110111011001100110;
rgb[7526] = 24'b001111011000111001111011;
rgb[7527] = 24'b010001111010011010001111;
rgb[7528] = 24'b010110001011011110100000;
rgb[7529] = 24'b011100001100000110101110;
rgb[7530] = 24'b100001111100110010111011;
rgb[7531] = 24'b100111111101011011001001;
rgb[7532] = 24'b101101111110000011010110;
rgb[7533] = 24'b110011111110101011100100;
rgb[7534] = 24'b111001111111010011110001;
rgb[7535] = 24'b111111111111111011111110;
rgb[7536] = 24'b000000000000000000000000;
rgb[7537] = 24'b000010010001100000010101;
rgb[7538] = 24'b000100100011000100101010;
rgb[7539] = 24'b000110110100101000111111;
rgb[7540] = 24'b001001000110001101010100;
rgb[7541] = 24'b001011010111110001101001;
rgb[7542] = 24'b001101101001010101111110;
rgb[7543] = 24'b001111111010111010010100;
rgb[7544] = 24'b010100001011111110100101;
rgb[7545] = 24'b011010011100100010110001;
rgb[7546] = 24'b100000101101000110111110;
rgb[7547] = 24'b100110111101101011001011;
rgb[7548] = 24'b101101001110001111011000;
rgb[7549] = 24'b110011011110110011100101;
rgb[7550] = 24'b111001101111010111110010;
rgb[7551] = 24'b111111111111111111111111;
rgb[7552] = 24'b000000000000000000000000;
rgb[7553] = 24'b000001110001101000010101;
rgb[7554] = 24'b000011110011010000101011;
rgb[7555] = 24'b000101110100111001000001;
rgb[7556] = 24'b000111110110100001010110;
rgb[7557] = 24'b001001111000001001101100;
rgb[7558] = 24'b001011111001110010000010;
rgb[7559] = 24'b001101111011011010011000;
rgb[7560] = 24'b010010001100011110101001;
rgb[7561] = 24'b011000101100111110110101;
rgb[7562] = 24'b011111001101011111000001;
rgb[7563] = 24'b100101101101111111001101;
rgb[7564] = 24'b101100001110011111011010;
rgb[7565] = 24'b110010101110111111100110;
rgb[7566] = 24'b111001001111011111110010;
rgb[7567] = 24'b111111111111111011111110;
rgb[7568] = 24'b000000000000000000000000;
rgb[7569] = 24'b000001100001101100010110;
rgb[7570] = 24'b000011010011011000101100;
rgb[7571] = 24'b000101000101000101000011;
rgb[7572] = 24'b000110110110110001011001;
rgb[7573] = 24'b001000011000100001101111;
rgb[7574] = 24'b001010001010001110000110;
rgb[7575] = 24'b001011111011111010011100;
rgb[7576] = 24'b010000001100111110101101;
rgb[7577] = 24'b010110111101011010111001;
rgb[7578] = 24'b011101101101110111000100;
rgb[7579] = 24'b100100101110001111010000;
rgb[7580] = 24'b101011011110101011011100;
rgb[7581] = 24'b110010001111000111100111;
rgb[7582] = 24'b111000111111100011110011;
rgb[7583] = 24'b111111111111111111111111;
rgb[7584] = 24'b000000000000000000000000;
rgb[7585] = 24'b000001010001110000010110;
rgb[7586] = 24'b000010110011100000101101;
rgb[7587] = 24'b000100010101010101000100;
rgb[7588] = 24'b000101100111000101011011;
rgb[7589] = 24'b000111001000110101110010;
rgb[7590] = 24'b001000101010101010001001;
rgb[7591] = 24'b001001111100011010100000;
rgb[7592] = 24'b001110001101011110110001;
rgb[7593] = 24'b010101001101110110111100;
rgb[7594] = 24'b011100011110001011000111;
rgb[7595] = 24'b100011011110100011010010;
rgb[7596] = 24'b101010101110111011011101;
rgb[7597] = 24'b110001101111001111101000;
rgb[7598] = 24'b111000101111100111110011;
rgb[7599] = 24'b111111111111111011111110;
rgb[7600] = 24'b000000000000000000000000;
rgb[7601] = 24'b000001000001110100010111;
rgb[7602] = 24'b000010010011101000101111;
rgb[7603] = 24'b000011010101100001000110;
rgb[7604] = 24'b000100100111010101011110;
rgb[7605] = 24'b000101101001001101110101;
rgb[7606] = 24'b000110111011000010001101;
rgb[7607] = 24'b000111111100111010100100;
rgb[7608] = 24'b001100001101111110110101;
rgb[7609] = 24'b010011101110001111000000;
rgb[7610] = 24'b011010111110100011001010;
rgb[7611] = 24'b100010011110110011010101;
rgb[7612] = 24'b101001101111000111011111;
rgb[7613] = 24'b110001001111010111101010;
rgb[7614] = 24'b111000011111101011110100;
rgb[7615] = 24'b111111111111111111111111;
rgb[7616] = 24'b000000000000000000000000;
rgb[7617] = 24'b000000110001111000011000;
rgb[7618] = 24'b000001100011110100110000;
rgb[7619] = 24'b000010100101101101001000;
rgb[7620] = 24'b000011010111101001100000;
rgb[7621] = 24'b000100001001100101111000;
rgb[7622] = 24'b000101001011011110010000;
rgb[7623] = 24'b000101111101011010101000;
rgb[7624] = 24'b001010001110011110111001;
rgb[7625] = 24'b010001111110101011000011;
rgb[7626] = 24'b011001011110111011001101;
rgb[7627] = 24'b100001001111000111010111;
rgb[7628] = 24'b101000111111010011100001;
rgb[7629] = 24'b110000011111100011101011;
rgb[7630] = 24'b111000001111101111110101;
rgb[7631] = 24'b111111111111111111111111;
rgb[7632] = 24'b000000000000000000000000;
rgb[7633] = 24'b000000100001111100011000;
rgb[7634] = 24'b000001000011111100110001;
rgb[7635] = 24'b000001100101111101001010;
rgb[7636] = 24'b000010010111111001100010;
rgb[7637] = 24'b000010111001111001111011;
rgb[7638] = 24'b000011011011111010010100;
rgb[7639] = 24'b000011111101111010101101;
rgb[7640] = 24'b001000001110111110111110;
rgb[7641] = 24'b010000001111000111000111;
rgb[7642] = 24'b011000001111001111010000;
rgb[7643] = 24'b100000001111010111011001;
rgb[7644] = 24'b100111111111100011100011;
rgb[7645] = 24'b101111111111101011101100;
rgb[7646] = 24'b110111111111110011110101;
rgb[7647] = 24'b111111111111111111111111;
rgb[7648] = 24'b000000000000000000000000;
rgb[7649] = 24'b000000010010000000011001;
rgb[7650] = 24'b000000100100000100110010;
rgb[7651] = 24'b000000110110001001001011;
rgb[7652] = 24'b000001001000001101100101;
rgb[7653] = 24'b000001011010010001111110;
rgb[7654] = 24'b000001101100010110010111;
rgb[7655] = 24'b000001111110011010110001;
rgb[7656] = 24'b000110001111011111000010;
rgb[7657] = 24'b001110011111100011001010;
rgb[7658] = 24'b010110101111100111010011;
rgb[7659] = 24'b011110111111101011011100;
rgb[7660] = 24'b100111001111101111100100;
rgb[7661] = 24'b101111011111110011101101;
rgb[7662] = 24'b110111101111110111110110;
rgb[7663] = 24'b111111111111111111111111;
rgb[7664] = 24'b000000000000000000000000;
rgb[7665] = 24'b000000000010001000011001;
rgb[7666] = 24'b000000000100010000110011;
rgb[7667] = 24'b000000000110011001001101;
rgb[7668] = 24'b000000001000100001100111;
rgb[7669] = 24'b000000001010101010000001;
rgb[7670] = 24'b000000001100110010011011;
rgb[7671] = 24'b000000001110111010110101;
rgb[7672] = 24'b000100011111111011000110;
rgb[7673] = 24'b001100101111111111001110;
rgb[7674] = 24'b010101011111111011010110;
rgb[7675] = 24'b011101101111111111011110;
rgb[7676] = 24'b100110011111111111100110;
rgb[7677] = 24'b101110111111111111101110;
rgb[7678] = 24'b110111011111111111110110;
rgb[7679] = 24'b111111111111111111111111;
rgb[7680] = 24'b000000000000000000000000;
rgb[7681] = 24'b000100010001000100010001;
rgb[7682] = 24'b001000100010001000100010;
rgb[7683] = 24'b001100110011001100110011;
rgb[7684] = 24'b010001000100010001000100;
rgb[7685] = 24'b010101010101010101010101;
rgb[7686] = 24'b011001100110011001100110;
rgb[7687] = 24'b011101110111011101110111;
rgb[7688] = 24'b100010001000100010001000;
rgb[7689] = 24'b100110011001100110011001;
rgb[7690] = 24'b101010101010101010101010;
rgb[7691] = 24'b101110111011101110111011;
rgb[7692] = 24'b110011001100110011001100;
rgb[7693] = 24'b110111011101110111011101;
rgb[7694] = 24'b111011101110111011101110;
rgb[7695] = 24'b111111111111111111111111;
rgb[7696] = 24'b000000000000000000000000;
rgb[7697] = 24'b000011110001001000010001;
rgb[7698] = 24'b000111110010010000100011;
rgb[7699] = 24'b001011110011011000110101;
rgb[7700] = 24'b001111110100100001000111;
rgb[7701] = 24'b010011110101101001011001;
rgb[7702] = 24'b010111110110110001101010;
rgb[7703] = 24'b011011110111111001111100;
rgb[7704] = 24'b100000001000111110001101;
rgb[7705] = 24'b100100101001111110011101;
rgb[7706] = 24'b101001001010111110101110;
rgb[7707] = 24'b101101101011111110111110;
rgb[7708] = 24'b110010001100111111001110;
rgb[7709] = 24'b110110101101111111011110;
rgb[7710] = 24'b111011001110111111101110;
rgb[7711] = 24'b111111111111111111111111;
rgb[7712] = 24'b000000000000000000000000;
rgb[7713] = 24'b000011100001001100010010;
rgb[7714] = 24'b000111010010011000100101;
rgb[7715] = 24'b001011000011100100110111;
rgb[7716] = 24'b001110100100110101001010;
rgb[7717] = 24'b010010010110000001011101;
rgb[7718] = 24'b010110000111001101101111;
rgb[7719] = 24'b011001111000011010000010;
rgb[7720] = 24'b011110001001011110010011;
rgb[7721] = 24'b100010111010011010100010;
rgb[7722] = 24'b100111101011010110110010;
rgb[7723] = 24'b101100011100010011000001;
rgb[7724] = 24'b110001011101001011010000;
rgb[7725] = 24'b110110001110000111100000;
rgb[7726] = 24'b111010111111000011101111;
rgb[7727] = 24'b111111111111111111111111;
rgb[7728] = 24'b000000000000000000000000;
rgb[7729] = 24'b000011010001010000010011;
rgb[7730] = 24'b000110110010100000100110;
rgb[7731] = 24'b001010000011110100111010;
rgb[7732] = 24'b001101100101000101001101;
rgb[7733] = 24'b010001000110010101100001;
rgb[7734] = 24'b010100010111101001110100;
rgb[7735] = 24'b010111111000111010001000;
rgb[7736] = 24'b011100001001111110011001;
rgb[7737] = 24'b100001001010110110100111;
rgb[7738] = 24'b100110001011101110110110;
rgb[7739] = 24'b101011011100100011000100;
rgb[7740] = 24'b110000011101011011010011;
rgb[7741] = 24'b110101101110001111100001;
rgb[7742] = 24'b111010101111000111110000;
rgb[7743] = 24'b111111111111111111111111;
rgb[7744] = 24'b000000000000000000000000;
rgb[7745] = 24'b000011000001010100010100;
rgb[7746] = 24'b000110000010101100101000;
rgb[7747] = 24'b001001010100000000111100;
rgb[7748] = 24'b001100010101011001010000;
rgb[7749] = 24'b001111100110101101100101;
rgb[7750] = 24'b010010101000000101111001;
rgb[7751] = 24'b010101111001011010001101;
rgb[7752] = 24'b011010001010011110011110;
rgb[7753] = 24'b011111011011010010101100;
rgb[7754] = 24'b100100111100000010111010;
rgb[7755] = 24'b101010001100110111000111;
rgb[7756] = 24'b101111101101100111010101;
rgb[7757] = 24'b110100111110011011100011;
rgb[7758] = 24'b111010011111001011110001;
rgb[7759] = 24'b111111111111111111111111;
rgb[7760] = 24'b000000000000000000000000;
rgb[7761] = 24'b000010110001011000010101;
rgb[7762] = 24'b000101100010110100101010;
rgb[7763] = 24'b001000100100010000111111;
rgb[7764] = 24'b001011010101101001010100;
rgb[7765] = 24'b001110000111000101101001;
rgb[7766] = 24'b010001001000100001111110;
rgb[7767] = 24'b010011111001111010010011;
rgb[7768] = 24'b011000001010111110100100;
rgb[7769] = 24'b011101101011101110110001;
rgb[7770] = 24'b100011011100011010111110;
rgb[7771] = 24'b101001001101000111001011;
rgb[7772] = 24'b101110111101110111011000;
rgb[7773] = 24'b110100011110100011100101;
rgb[7774] = 24'b111010001111001111110010;
rgb[7775] = 24'b111111111111111111111111;
rgb[7776] = 24'b000000000000000000000000;
rgb[7777] = 24'b000010100001011100010101;
rgb[7778] = 24'b000101000010111100101011;
rgb[7779] = 24'b000111100100011101000001;
rgb[7780] = 24'b001010000101111101010111;
rgb[7781] = 24'b001100110111011001101101;
rgb[7782] = 24'b001111011000111010000011;
rgb[7783] = 24'b010001111010011010011001;
rgb[7784] = 24'b010110001011011110101010;
rgb[7785] = 24'b011100001100000110110110;
rgb[7786] = 24'b100001111100110011000010;
rgb[7787] = 24'b100111111101011011001110;
rgb[7788] = 24'b101101111110000011011010;
rgb[7789] = 24'b110011111110101011100110;
rgb[7790] = 24'b111001111111010011110010;
rgb[7791] = 24'b111111111111111011111110;
rgb[7792] = 24'b000000000000000000000000;
rgb[7793] = 24'b000010010001100000010110;
rgb[7794] = 24'b000100100011000100101101;
rgb[7795] = 24'b000110110100101001000100;
rgb[7796] = 24'b001001000110001101011010;
rgb[7797] = 24'b001011010111110001110001;
rgb[7798] = 24'b001101101001010110001000;
rgb[7799] = 24'b001111111010111010011110;
rgb[7800] = 24'b010100001011111110101111;
rgb[7801] = 24'b011010011100100010111011;
rgb[7802] = 24'b100000101101000111000110;
rgb[7803] = 24'b100110111101101011010001;
rgb[7804] = 24'b101101001110001111011101;
rgb[7805] = 24'b110011011110110011101000;
rgb[7806] = 24'b111001101111010111110011;
rgb[7807] = 24'b111111111111111111111111;
rgb[7808] = 24'b000000000000000000000000;
rgb[7809] = 24'b000001110001101000010111;
rgb[7810] = 24'b000011110011010000101110;
rgb[7811] = 24'b000101110100111001000110;
rgb[7812] = 24'b000111110110100001011101;
rgb[7813] = 24'b001001111000001001110101;
rgb[7814] = 24'b001011111001110010001100;
rgb[7815] = 24'b001101111011011010100100;
rgb[7816] = 24'b010010001100011110110101;
rgb[7817] = 24'b011000101100111110111111;
rgb[7818] = 24'b011111001101011111001010;
rgb[7819] = 24'b100101101101111111010100;
rgb[7820] = 24'b101100001110011111011111;
rgb[7821] = 24'b110010101110111111101001;
rgb[7822] = 24'b111001001111011111110100;
rgb[7823] = 24'b111111111111111011111110;
rgb[7824] = 24'b000000000000000000000000;
rgb[7825] = 24'b000001100001101100011000;
rgb[7826] = 24'b000011010011011000110000;
rgb[7827] = 24'b000101000101000101001000;
rgb[7828] = 24'b000110110110110001100001;
rgb[7829] = 24'b001000011000100001111001;
rgb[7830] = 24'b001010001010001110010001;
rgb[7831] = 24'b001011111011111010101010;
rgb[7832] = 24'b010000001100111110111011;
rgb[7833] = 24'b010110111101011011000100;
rgb[7834] = 24'b011101101101110111001110;
rgb[7835] = 24'b100100101110001111011000;
rgb[7836] = 24'b101011011110101011100001;
rgb[7837] = 24'b110010001111000111101011;
rgb[7838] = 24'b111000111111100011110101;
rgb[7839] = 24'b111111111111111111111111;
rgb[7840] = 24'b000000000000000000000000;
rgb[7841] = 24'b000001010001110000011001;
rgb[7842] = 24'b000010110011100000110010;
rgb[7843] = 24'b000100010101010101001011;
rgb[7844] = 24'b000101100111000101100100;
rgb[7845] = 24'b000111001000110101111101;
rgb[7846] = 24'b001000101010101010010110;
rgb[7847] = 24'b001001111100011010101111;
rgb[7848] = 24'b001110001101011111000000;
rgb[7849] = 24'b010101001101110111001001;
rgb[7850] = 24'b011100011110001011010010;
rgb[7851] = 24'b100011011110100011011011;
rgb[7852] = 24'b101010101110111011100100;
rgb[7853] = 24'b110001101111001111101101;
rgb[7854] = 24'b111000101111100111110110;
rgb[7855] = 24'b111111111111111011111110;
rgb[7856] = 24'b000000000000000000000000;
rgb[7857] = 24'b000001000001110100011001;
rgb[7858] = 24'b000010010011101000110011;
rgb[7859] = 24'b000011010101100001001101;
rgb[7860] = 24'b000100100111010101100111;
rgb[7861] = 24'b000101101001001110000001;
rgb[7862] = 24'b000110111011000010011011;
rgb[7863] = 24'b000111111100111010110101;
rgb[7864] = 24'b001100001101111111000110;
rgb[7865] = 24'b010011101110001111001110;
rgb[7866] = 24'b011010111110100011010110;
rgb[7867] = 24'b100010011110110011011110;
rgb[7868] = 24'b101001101111000111100110;
rgb[7869] = 24'b110001001111010111101110;
rgb[7870] = 24'b111000011111101011110110;
rgb[7871] = 24'b111111111111111111111111;
rgb[7872] = 24'b000000000000000000000000;
rgb[7873] = 24'b000000110001111000011010;
rgb[7874] = 24'b000001100011110100110101;
rgb[7875] = 24'b000010100101101101010000;
rgb[7876] = 24'b000011010111101001101010;
rgb[7877] = 24'b000100001001100110000101;
rgb[7878] = 24'b000101001011011110100000;
rgb[7879] = 24'b000101111101011010111011;
rgb[7880] = 24'b001010001110011111001100;
rgb[7881] = 24'b010001111110101011010011;
rgb[7882] = 24'b011001011110111011011010;
rgb[7883] = 24'b100001001111000111100001;
rgb[7884] = 24'b101000111111010011101001;
rgb[7885] = 24'b110000011111100011110000;
rgb[7886] = 24'b111000001111101111110111;
rgb[7887] = 24'b111111111111111111111111;
rgb[7888] = 24'b000000000000000000000000;
rgb[7889] = 24'b000000100001111100011011;
rgb[7890] = 24'b000001000011111100110111;
rgb[7891] = 24'b000001100101111101010010;
rgb[7892] = 24'b000010010111111001101110;
rgb[7893] = 24'b000010111001111010001001;
rgb[7894] = 24'b000011011011111010100101;
rgb[7895] = 24'b000011111101111011000000;
rgb[7896] = 24'b001000001110111111010001;
rgb[7897] = 24'b010000001111000111011000;
rgb[7898] = 24'b011000001111001111011110;
rgb[7899] = 24'b100000001111010111100101;
rgb[7900] = 24'b100111111111100011101011;
rgb[7901] = 24'b101111111111101011110010;
rgb[7902] = 24'b110111111111110011111000;
rgb[7903] = 24'b111111111111111111111111;
rgb[7904] = 24'b000000000000000000000000;
rgb[7905] = 24'b000000010010000000011100;
rgb[7906] = 24'b000000100100000100111000;
rgb[7907] = 24'b000000110110001001010101;
rgb[7908] = 24'b000001001000001101110001;
rgb[7909] = 24'b000001011010010010001101;
rgb[7910] = 24'b000001101100010110101010;
rgb[7911] = 24'b000001111110011011000110;
rgb[7912] = 24'b000110001111011111010111;
rgb[7913] = 24'b001110011111100011011100;
rgb[7914] = 24'b010110101111100111100010;
rgb[7915] = 24'b011110111111101011101000;
rgb[7916] = 24'b100111001111101111101110;
rgb[7917] = 24'b101111011111110011110011;
rgb[7918] = 24'b110111101111110111111001;
rgb[7919] = 24'b111111111111111111111111;
rgb[7920] = 24'b000000000000000000000000;
rgb[7921] = 24'b000000000010001000011101;
rgb[7922] = 24'b000000000100010000111010;
rgb[7923] = 24'b000000000110011001010111;
rgb[7924] = 24'b000000001000100001110100;
rgb[7925] = 24'b000000001010101010010001;
rgb[7926] = 24'b000000001100110010101110;
rgb[7927] = 24'b000000001110111011001100;
rgb[7928] = 24'b000100011111111011011100;
rgb[7929] = 24'b001100101111111111100001;
rgb[7930] = 24'b010101011111111011100110;
rgb[7931] = 24'b011101101111111111101011;
rgb[7932] = 24'b100110011111111111110000;
rgb[7933] = 24'b101110111111111111110101;
rgb[7934] = 24'b110111011111111111111010;
rgb[7935] = 24'b111111111111111111111111;
rgb[7936] = 24'b000000000000000000000000;
rgb[7937] = 24'b000100010001000100010001;
rgb[7938] = 24'b001000100010001000100010;
rgb[7939] = 24'b001100110011001100110011;
rgb[7940] = 24'b010001000100010001000100;
rgb[7941] = 24'b010101010101010101010101;
rgb[7942] = 24'b011001100110011001100110;
rgb[7943] = 24'b011101110111011101110111;
rgb[7944] = 24'b100010001000100010001000;
rgb[7945] = 24'b100110011001100110011001;
rgb[7946] = 24'b101010101010101010101010;
rgb[7947] = 24'b101110111011101110111011;
rgb[7948] = 24'b110011001100110011001100;
rgb[7949] = 24'b110111011101110111011101;
rgb[7950] = 24'b111011101110111011101110;
rgb[7951] = 24'b111111111111111111111111;
rgb[7952] = 24'b000000000000000000000000;
rgb[7953] = 24'b000011110001001000010010;
rgb[7954] = 24'b000111110010010000100100;
rgb[7955] = 24'b001011110011011000110110;
rgb[7956] = 24'b001111110100100001001000;
rgb[7957] = 24'b010011110101101001011010;
rgb[7958] = 24'b010111110110110001101100;
rgb[7959] = 24'b011011110111111001111110;
rgb[7960] = 24'b100000001000111110001111;
rgb[7961] = 24'b100100101001111110011111;
rgb[7962] = 24'b101001001010111110101111;
rgb[7963] = 24'b101101101011111110111111;
rgb[7964] = 24'b110010001100111111001111;
rgb[7965] = 24'b110110101101111111011111;
rgb[7966] = 24'b111011001110111111101111;
rgb[7967] = 24'b111111111111111111111111;
rgb[7968] = 24'b000000000000000000000000;
rgb[7969] = 24'b000011100001001100010011;
rgb[7970] = 24'b000111010010011000100110;
rgb[7971] = 24'b001011000011100100111001;
rgb[7972] = 24'b001110100100110101001100;
rgb[7973] = 24'b010010010110000001011111;
rgb[7974] = 24'b010110000111001101110010;
rgb[7975] = 24'b011001111000011010000101;
rgb[7976] = 24'b011110001001011110010110;
rgb[7977] = 24'b100010111010011010100101;
rgb[7978] = 24'b100111101011010110110100;
rgb[7979] = 24'b101100011100010011000011;
rgb[7980] = 24'b110001011101001011010010;
rgb[7981] = 24'b110110001110000111100001;
rgb[7982] = 24'b111010111111000011110000;
rgb[7983] = 24'b111111111111111111111111;
rgb[7984] = 24'b000000000000000000000000;
rgb[7985] = 24'b000011010001010000010100;
rgb[7986] = 24'b000110110010100000101000;
rgb[7987] = 24'b001010000011110100111100;
rgb[7988] = 24'b001101100101000101010000;
rgb[7989] = 24'b010001000110010101100100;
rgb[7990] = 24'b010100010111101001111000;
rgb[7991] = 24'b010111111000111010001100;
rgb[7992] = 24'b011100001001111110011101;
rgb[7993] = 24'b100001001010110110101011;
rgb[7994] = 24'b100110001011101110111001;
rgb[7995] = 24'b101011011100100011000111;
rgb[7996] = 24'b110000011101011011010101;
rgb[7997] = 24'b110101101110001111100011;
rgb[7998] = 24'b111010101111000111110001;
rgb[7999] = 24'b111111111111111111111111;
rgb[8000] = 24'b000000000000000000000000;
rgb[8001] = 24'b000011000001010100010101;
rgb[8002] = 24'b000110000010101100101010;
rgb[8003] = 24'b001001010100000000111111;
rgb[8004] = 24'b001100010101011001010100;
rgb[8005] = 24'b001111100110101101101001;
rgb[8006] = 24'b010010101000000101111110;
rgb[8007] = 24'b010101111001011010010011;
rgb[8008] = 24'b011010001010011110100100;
rgb[8009] = 24'b011111011011010010110001;
rgb[8010] = 24'b100100111100000010111110;
rgb[8011] = 24'b101010001100110111001011;
rgb[8012] = 24'b101111101101100111011000;
rgb[8013] = 24'b110100111110011011100101;
rgb[8014] = 24'b111010011111001011110010;
rgb[8015] = 24'b111111111111111111111111;
rgb[8016] = 24'b000000000000000000000000;
rgb[8017] = 24'b000010110001011000010110;
rgb[8018] = 24'b000101100010110100101100;
rgb[8019] = 24'b001000100100010001000010;
rgb[8020] = 24'b001011010101101001011000;
rgb[8021] = 24'b001110000111000101101110;
rgb[8022] = 24'b010001001000100010000100;
rgb[8023] = 24'b010011111001111010011010;
rgb[8024] = 24'b011000001010111110101011;
rgb[8025] = 24'b011101101011101110110111;
rgb[8026] = 24'b100011011100011011000011;
rgb[8027] = 24'b101001001101000111001111;
rgb[8028] = 24'b101110111101110111011011;
rgb[8029] = 24'b110100011110100011100111;
rgb[8030] = 24'b111010001111001111110011;
rgb[8031] = 24'b111111111111111111111111;
rgb[8032] = 24'b000000000000000000000000;
rgb[8033] = 24'b000010100001011100010111;
rgb[8034] = 24'b000101000010111100101110;
rgb[8035] = 24'b000111100100011101000101;
rgb[8036] = 24'b001010000101111101011100;
rgb[8037] = 24'b001100110111011001110011;
rgb[8038] = 24'b001111011000111010001010;
rgb[8039] = 24'b010001111010011010100010;
rgb[8040] = 24'b010110001011011110110011;
rgb[8041] = 24'b011100001100000110111101;
rgb[8042] = 24'b100001111100110011001000;
rgb[8043] = 24'b100111111101011011010011;
rgb[8044] = 24'b101101111110000011011110;
rgb[8045] = 24'b110011111110101011101001;
rgb[8046] = 24'b111001111111010011110100;
rgb[8047] = 24'b111111111111111011111110;
rgb[8048] = 24'b000000000000000000000000;
rgb[8049] = 24'b000010010001100000011000;
rgb[8050] = 24'b000100100011000100110000;
rgb[8051] = 24'b000110110100101001001000;
rgb[8052] = 24'b001001000110001101100000;
rgb[8053] = 24'b001011010111110001111000;
rgb[8054] = 24'b001101101001010110010001;
rgb[8055] = 24'b001111111010111010101001;
rgb[8056] = 24'b010100001011111110111010;
rgb[8057] = 24'b011010011100100011000100;
rgb[8058] = 24'b100000101101000111001101;
rgb[8059] = 24'b100110111101101011010111;
rgb[8060] = 24'b101101001110001111100001;
rgb[8061] = 24'b110011011110110011101011;
rgb[8062] = 24'b111001101111010111110101;
rgb[8063] = 24'b111111111111111111111111;
rgb[8064] = 24'b000000000000000000000000;
rgb[8065] = 24'b000001110001101000011001;
rgb[8066] = 24'b000011110011010000110010;
rgb[8067] = 24'b000101110100111001001011;
rgb[8068] = 24'b000111110110100001100100;
rgb[8069] = 24'b001001111000001001111110;
rgb[8070] = 24'b001011111001110010010111;
rgb[8071] = 24'b001101111011011010110000;
rgb[8072] = 24'b010010001100011111000001;
rgb[8073] = 24'b011000101100111111001010;
rgb[8074] = 24'b011111001101011111010011;
rgb[8075] = 24'b100101101101111111011011;
rgb[8076] = 24'b101100001110011111100100;
rgb[8077] = 24'b110010101110111111101101;
rgb[8078] = 24'b111001001111011111110110;
rgb[8079] = 24'b111111111111111011111110;
rgb[8080] = 24'b000000000000000000000000;
rgb[8081] = 24'b000001100001101100011010;
rgb[8082] = 24'b000011010011011000110100;
rgb[8083] = 24'b000101000101000101001110;
rgb[8084] = 24'b000110110110110001101000;
rgb[8085] = 24'b001000011000100010000011;
rgb[8086] = 24'b001010001010001110011101;
rgb[8087] = 24'b001011111011111010110111;
rgb[8088] = 24'b010000001100111111001000;
rgb[8089] = 24'b010110111101011011010000;
rgb[8090] = 24'b011101101101110111011000;
rgb[8091] = 24'b100100101110001111011111;
rgb[8092] = 24'b101011011110101011100111;
rgb[8093] = 24'b110010001111000111101111;
rgb[8094] = 24'b111000111111100011110111;
rgb[8095] = 24'b111111111111111111111111;
rgb[8096] = 24'b000000000000000000000000;
rgb[8097] = 24'b000001010001110000011011;
rgb[8098] = 24'b000010110011100000110110;
rgb[8099] = 24'b000100010101010101010001;
rgb[8100] = 24'b000101100111000101101101;
rgb[8101] = 24'b000111001000110110001000;
rgb[8102] = 24'b001000101010101010100011;
rgb[8103] = 24'b001001111100011010111110;
rgb[8104] = 24'b001110001101011111001111;
rgb[8105] = 24'b010101001101110111010110;
rgb[8106] = 24'b011100011110001011011101;
rgb[8107] = 24'b100011011110100011100100;
rgb[8108] = 24'b101010101110111011101010;
rgb[8109] = 24'b110001101111001111110001;
rgb[8110] = 24'b111000101111100111111000;
rgb[8111] = 24'b111111111111111011111110;
rgb[8112] = 24'b000000000000000000000000;
rgb[8113] = 24'b000001000001110100011100;
rgb[8114] = 24'b000010010011101000111000;
rgb[8115] = 24'b000011010101100001010100;
rgb[8116] = 24'b000100100111010101110001;
rgb[8117] = 24'b000101101001001110001101;
rgb[8118] = 24'b000110111011000010101001;
rgb[8119] = 24'b000111111100111011000101;
rgb[8120] = 24'b001100001101111111010110;
rgb[8121] = 24'b010011101110001111011100;
rgb[8122] = 24'b011010111110100011100010;
rgb[8123] = 24'b100010011110110011101000;
rgb[8124] = 24'b101001101111000111101101;
rgb[8125] = 24'b110001001111010111110011;
rgb[8126] = 24'b111000011111101011111001;
rgb[8127] = 24'b111111111111111111111111;
rgb[8128] = 24'b000000000000000000000000;
rgb[8129] = 24'b000000110001111000011101;
rgb[8130] = 24'b000001100011110100111010;
rgb[8131] = 24'b000010100101101101010111;
rgb[8132] = 24'b000011010111101001110101;
rgb[8133] = 24'b000100001001100110010010;
rgb[8134] = 24'b000101001011011110101111;
rgb[8135] = 24'b000101111101011011001101;
rgb[8136] = 24'b001010001110011111011110;
rgb[8137] = 24'b010001111110101011100010;
rgb[8138] = 24'b011001011110111011100111;
rgb[8139] = 24'b100001001111000111101100;
rgb[8140] = 24'b101000111111010011110000;
rgb[8141] = 24'b110000011111100011110101;
rgb[8142] = 24'b111000001111101111111010;
rgb[8143] = 24'b111111111111111111111111;
rgb[8144] = 24'b000000000000000000000000;
rgb[8145] = 24'b000000100001111100011110;
rgb[8146] = 24'b000001000011111100111100;
rgb[8147] = 24'b000001100101111101011010;
rgb[8148] = 24'b000010010111111001111001;
rgb[8149] = 24'b000010111001111010010111;
rgb[8150] = 24'b000011011011111010110101;
rgb[8151] = 24'b000011111101111011010100;
rgb[8152] = 24'b001000001110111111100101;
rgb[8153] = 24'b010000001111000111101000;
rgb[8154] = 24'b011000001111001111101100;
rgb[8155] = 24'b100000001111010111110000;
rgb[8156] = 24'b100111111111100011110011;
rgb[8157] = 24'b101111111111101011110111;
rgb[8158] = 24'b110111111111110011111011;
rgb[8159] = 24'b111111111111111111111111;
rgb[8160] = 24'b000000000000000000000000;
rgb[8161] = 24'b000000010010000000011111;
rgb[8162] = 24'b000000100100000100111110;
rgb[8163] = 24'b000000110110001001011110;
rgb[8164] = 24'b000001001000001101111101;
rgb[8165] = 24'b000001011010010010011100;
rgb[8166] = 24'b000001101100010110111100;
rgb[8167] = 24'b000001111110011011011011;
rgb[8168] = 24'b000110001111011111101100;
rgb[8169] = 24'b001110011111100011101111;
rgb[8170] = 24'b010110101111100111110001;
rgb[8171] = 24'b011110111111101011110100;
rgb[8172] = 24'b100111001111101111110111;
rgb[8173] = 24'b101111011111110011111001;
rgb[8174] = 24'b110111101111110111111100;
rgb[8175] = 24'b111111111111111111111111;
rgb[8176] = 24'b000000000000000000000000;
rgb[8177] = 24'b000000000010001000100000;
rgb[8178] = 24'b000000000100010001000000;
rgb[8179] = 24'b000000000110011001100001;
rgb[8180] = 24'b000000001000100010000001;
rgb[8181] = 24'b000000001010101010100001;
rgb[8182] = 24'b000000001100110011000010;
rgb[8183] = 24'b000000001110111011100010;
rgb[8184] = 24'b000100011111111011110011;
rgb[8185] = 24'b001100101111111111110101;
rgb[8186] = 24'b010101011111111011110110;
rgb[8187] = 24'b011101101111111111111000;
rgb[8188] = 24'b100110011111111111111010;
rgb[8189] = 24'b101110111111111111111011;
rgb[8190] = 24'b110111011111111111111101;
rgb[8191] = 24'b111111111111111111111111;
rgb[8192] = 24'b000000000000000000000000;
rgb[8193] = 24'b000100010001000100010001;
rgb[8194] = 24'b001000100010001000100010;
rgb[8195] = 24'b001100110011001100110011;
rgb[8196] = 24'b010001000100010001000100;
rgb[8197] = 24'b010101010101010101010101;
rgb[8198] = 24'b011001100110011001100110;
rgb[8199] = 24'b011101110111011101110111;
rgb[8200] = 24'b100010001000100010001000;
rgb[8201] = 24'b100110011001100110011001;
rgb[8202] = 24'b101010101010101010101010;
rgb[8203] = 24'b101110111011101110111011;
rgb[8204] = 24'b110011001100110011001100;
rgb[8205] = 24'b110111011101110111011101;
rgb[8206] = 24'b111011101110111011101110;
rgb[8207] = 24'b111111111111111111111111;
rgb[8208] = 24'b000000000000000000000000;
rgb[8209] = 24'b000011110001001000010010;
rgb[8210] = 24'b000111110010010000100100;
rgb[8211] = 24'b001011110011011000110110;
rgb[8212] = 24'b001111110100100001001000;
rgb[8213] = 24'b010011110101101001011010;
rgb[8214] = 24'b010111110110110001101100;
rgb[8215] = 24'b011011110111111001111110;
rgb[8216] = 24'b100000001000111110001111;
rgb[8217] = 24'b100100101001111110011111;
rgb[8218] = 24'b101001001010111110101111;
rgb[8219] = 24'b101101101011111110111111;
rgb[8220] = 24'b110010001100111111001111;
rgb[8221] = 24'b110110101101111111011111;
rgb[8222] = 24'b111011001110111111101111;
rgb[8223] = 24'b111111111111111111111111;
rgb[8224] = 24'b000000000000000000000000;
rgb[8225] = 24'b000011100001001100010011;
rgb[8226] = 24'b000111010010011000100110;
rgb[8227] = 24'b001011000011100100111001;
rgb[8228] = 24'b001110100100110001001101;
rgb[8229] = 24'b010010010101111101100000;
rgb[8230] = 24'b010110000111001001110011;
rgb[8231] = 24'b011001111000010110000110;
rgb[8232] = 24'b011110001001011010010111;
rgb[8233] = 24'b100010111010010110100110;
rgb[8234] = 24'b100111101011010010110101;
rgb[8235] = 24'b101100011100001111000100;
rgb[8236] = 24'b110001011101001011010010;
rgb[8237] = 24'b110110001110000111100001;
rgb[8238] = 24'b111010111111000011110000;
rgb[8239] = 24'b111111111111111111111111;
rgb[8240] = 24'b000000000000000000000000;
rgb[8241] = 24'b000011010001010000010100;
rgb[8242] = 24'b000110110010100000101000;
rgb[8243] = 24'b001010000011110000111101;
rgb[8244] = 24'b001101100101000001010001;
rgb[8245] = 24'b010001000110010001100101;
rgb[8246] = 24'b010100010111100001111010;
rgb[8247] = 24'b010111111000110010001110;
rgb[8248] = 24'b011100001001110110011111;
rgb[8249] = 24'b100001001010101110101101;
rgb[8250] = 24'b100110001011100110111011;
rgb[8251] = 24'b101011011100011111001000;
rgb[8252] = 24'b110000011101010111010110;
rgb[8253] = 24'b110101101110001111100011;
rgb[8254] = 24'b111010101111000111110001;
rgb[8255] = 24'b111111111111111111111111;
rgb[8256] = 24'b000000000000000000000000;
rgb[8257] = 24'b000011000001010100010101;
rgb[8258] = 24'b000110000010101000101011;
rgb[8259] = 24'b001001010011111101000000;
rgb[8260] = 24'b001100010101010001010110;
rgb[8261] = 24'b001111100110100101101011;
rgb[8262] = 24'b010010100111111010000001;
rgb[8263] = 24'b010101111001001110010110;
rgb[8264] = 24'b011010001010010010100111;
rgb[8265] = 24'b011111011011000110110100;
rgb[8266] = 24'b100100111011111011000000;
rgb[8267] = 24'b101010001100101111001101;
rgb[8268] = 24'b101111101101100011011001;
rgb[8269] = 24'b110100111110010111100110;
rgb[8270] = 24'b111010011111001011110010;
rgb[8271] = 24'b111111111111111111111111;
rgb[8272] = 24'b000000000000000000000000;
rgb[8273] = 24'b000010110001011000010110;
rgb[8274] = 24'b000101100010110000101101;
rgb[8275] = 24'b001000100100001001000100;
rgb[8276] = 24'b001011010101100001011010;
rgb[8277] = 24'b001110000110111001110001;
rgb[8278] = 24'b010001001000010010001000;
rgb[8279] = 24'b010011111001101010011110;
rgb[8280] = 24'b011000001010101110101111;
rgb[8281] = 24'b011101101011011110111011;
rgb[8282] = 24'b100011011100001111000110;
rgb[8283] = 24'b101001001100111111010001;
rgb[8284] = 24'b101110111101101111011101;
rgb[8285] = 24'b110100011110011111101000;
rgb[8286] = 24'b111010001111001111110011;
rgb[8287] = 24'b111111111111111111111111;
rgb[8288] = 24'b000000000000000000000000;
rgb[8289] = 24'b000010100001011100010111;
rgb[8290] = 24'b000101000010111000101111;
rgb[8291] = 24'b000111100100010101000111;
rgb[8292] = 24'b001010000101110001011111;
rgb[8293] = 24'b001100110111001101110110;
rgb[8294] = 24'b001111011000101010001110;
rgb[8295] = 24'b010001111010001010100110;
rgb[8296] = 24'b010110001011001110110111;
rgb[8297] = 24'b011100001011110111000001;
rgb[8298] = 24'b100001111100100011001100;
rgb[8299] = 24'b100111111101001111010110;
rgb[8300] = 24'b101101111101111011100000;
rgb[8301] = 24'b110011111110100111101010;
rgb[8302] = 24'b111001111111010011110100;
rgb[8303] = 24'b111111111111111011111110;
rgb[8304] = 24'b000000000000000000000000;
rgb[8305] = 24'b000010010001100000011000;
rgb[8306] = 24'b000100100011000000110001;
rgb[8307] = 24'b000110110100100001001010;
rgb[8308] = 24'b001001000110000001100011;
rgb[8309] = 24'b001011010111100001111100;
rgb[8310] = 24'b001101101001000110010101;
rgb[8311] = 24'b001111111010100110101110;
rgb[8312] = 24'b010100001011101010111111;
rgb[8313] = 24'b011010011100010011001000;
rgb[8314] = 24'b100000101100110111010001;
rgb[8315] = 24'b100110111101011111011010;
rgb[8316] = 24'b101101001110000111100011;
rgb[8317] = 24'b110011011110101111101100;
rgb[8318] = 24'b111001101111010111110101;
rgb[8319] = 24'b111111111111111111111111;
rgb[8320] = 24'b000000000000000000000000;
rgb[8321] = 24'b000001110001100100011010;
rgb[8322] = 24'b000011110011001000110100;
rgb[8323] = 24'b000101110100101101001110;
rgb[8324] = 24'b000111110110010001101000;
rgb[8325] = 24'b001001110111111010000010;
rgb[8326] = 24'b001011111001011110011100;
rgb[8327] = 24'b001101111011000010110110;
rgb[8328] = 24'b010010001100000111000111;
rgb[8329] = 24'b011000101100101011001111;
rgb[8330] = 24'b011111001101001111010111;
rgb[8331] = 24'b100101101101101111011111;
rgb[8332] = 24'b101100001110010011100111;
rgb[8333] = 24'b110010101110110111101111;
rgb[8334] = 24'b111001001111011011110111;
rgb[8335] = 24'b111111111111111011111110;
rgb[8336] = 24'b000000000000000000000000;
rgb[8337] = 24'b000001100001101000011011;
rgb[8338] = 24'b000011010011010000110110;
rgb[8339] = 24'b000101000100111001010001;
rgb[8340] = 24'b000110110110100001101100;
rgb[8341] = 24'b001000011000001110001000;
rgb[8342] = 24'b001010001001110110100011;
rgb[8343] = 24'b001011111011011110111110;
rgb[8344] = 24'b010000001100100011001111;
rgb[8345] = 24'b010110111101000011010110;
rgb[8346] = 24'b011101101101100011011101;
rgb[8347] = 24'b100100101101111111100011;
rgb[8348] = 24'b101011011110011111101010;
rgb[8349] = 24'b110010001110111111110001;
rgb[8350] = 24'b111000111111011111111000;
rgb[8351] = 24'b111111111111111111111111;
rgb[8352] = 24'b000000000000000000000000;
rgb[8353] = 24'b000001010001101100011100;
rgb[8354] = 24'b000010110011011000111000;
rgb[8355] = 24'b000100010101000101010101;
rgb[8356] = 24'b000101100110110101110001;
rgb[8357] = 24'b000111001000100010001101;
rgb[8358] = 24'b001000101010001110101010;
rgb[8359] = 24'b001001111011111011000110;
rgb[8360] = 24'b001110001100111111010111;
rgb[8361] = 24'b010101001101011011011101;
rgb[8362] = 24'b011100011101110111100010;
rgb[8363] = 24'b100011011110010011101000;
rgb[8364] = 24'b101010101110101011101110;
rgb[8365] = 24'b110001101111000111110011;
rgb[8366] = 24'b111000101111100011111001;
rgb[8367] = 24'b111111111111111011111110;
rgb[8368] = 24'b000000000000000000000000;
rgb[8369] = 24'b000001000001110000011101;
rgb[8370] = 24'b000010010011100000111010;
rgb[8371] = 24'b000011010101010001011000;
rgb[8372] = 24'b000100100111000101110101;
rgb[8373] = 24'b000101101000110110010011;
rgb[8374] = 24'b000110111010100110110000;
rgb[8375] = 24'b000111111100010111001110;
rgb[8376] = 24'b001100001101011011011111;
rgb[8377] = 24'b010011101101110011100011;
rgb[8378] = 24'b011010111110001011101000;
rgb[8379] = 24'b100010011110100011101100;
rgb[8380] = 24'b101001101110110111110001;
rgb[8381] = 24'b110001001111001111110101;
rgb[8382] = 24'b111000011111100111111010;
rgb[8383] = 24'b111111111111111111111111;
rgb[8384] = 24'b000000000000000000000000;
rgb[8385] = 24'b000000110001110100011110;
rgb[8386] = 24'b000001100011101000111101;
rgb[8387] = 24'b000010100101011101011011;
rgb[8388] = 24'b000011010111010101111010;
rgb[8389] = 24'b000100001001001010011001;
rgb[8390] = 24'b000101001010111110110111;
rgb[8391] = 24'b000101111100110111010110;
rgb[8392] = 24'b001010001101111011100111;
rgb[8393] = 24'b010001111110001011101010;
rgb[8394] = 24'b011001011110011111101110;
rgb[8395] = 24'b100001001110110011110001;
rgb[8396] = 24'b101000111111000011110100;
rgb[8397] = 24'b110000011111010111111000;
rgb[8398] = 24'b111000001111101011111011;
rgb[8399] = 24'b111111111111111111111111;
rgb[8400] = 24'b000000000000000000000000;
rgb[8401] = 24'b000000100001111000011111;
rgb[8402] = 24'b000001000011110000111111;
rgb[8403] = 24'b000001100101101001011111;
rgb[8404] = 24'b000010010111100101111110;
rgb[8405] = 24'b000010111001011110011110;
rgb[8406] = 24'b000011011011010110111110;
rgb[8407] = 24'b000011111101010011011110;
rgb[8408] = 24'b001000001110010111101111;
rgb[8409] = 24'b010000001110100011110001;
rgb[8410] = 24'b011000001110110011110011;
rgb[8411] = 24'b100000001111000011110101;
rgb[8412] = 24'b100111111111001111111000;
rgb[8413] = 24'b101111111111011111111010;
rgb[8414] = 24'b110111111111101111111100;
rgb[8415] = 24'b111111111111111111111111;
rgb[8416] = 24'b000000000000000000000000;
rgb[8417] = 24'b000000010001111100100000;
rgb[8418] = 24'b000000100011111001000001;
rgb[8419] = 24'b000000110101111001100010;
rgb[8420] = 24'b000001000111110110000011;
rgb[8421] = 24'b000001011001110010100100;
rgb[8422] = 24'b000001101011110011000101;
rgb[8423] = 24'b000001111101101111100110;
rgb[8424] = 24'b000110001110110011110111;
rgb[8425] = 24'b001110011110111111111000;
rgb[8426] = 24'b010110101111000111111001;
rgb[8427] = 24'b011110111111010011111010;
rgb[8428] = 24'b100111001111011111111011;
rgb[8429] = 24'b101111011111100111111100;
rgb[8430] = 24'b110111101111110011111101;
rgb[8431] = 24'b111111111111111111111111;
rgb[8432] = 24'b000000000000000000000000;
rgb[8433] = 24'b000000000010000000100010;
rgb[8434] = 24'b000000000100000001000100;
rgb[8435] = 24'b000000000110000101100110;
rgb[8436] = 24'b000000001000000110001000;
rgb[8437] = 24'b000000001010000110101010;
rgb[8438] = 24'b000000001100001011001100;
rgb[8439] = 24'b000000001110001011101110;
rgb[8440] = 24'b000100011111001111111110;
rgb[8441] = 24'b001100101111010111111111;
rgb[8442] = 24'b010101011111011011111110;
rgb[8443] = 24'b011101101111100011111111;
rgb[8444] = 24'b100110011111101011111111;
rgb[8445] = 24'b101110111111101111111111;
rgb[8446] = 24'b110111011111110111111111;
rgb[8447] = 24'b111111111111111111111111;
rgb[8448] = 24'b000000000000000000000000;
rgb[8449] = 24'b000100010001000100010001;
rgb[8450] = 24'b001000100010001000100010;
rgb[8451] = 24'b001100110011001100110011;
rgb[8452] = 24'b010001000100010001000100;
rgb[8453] = 24'b010101010101010101010101;
rgb[8454] = 24'b011001100110011001100110;
rgb[8455] = 24'b011101110111011101110111;
rgb[8456] = 24'b100010001000100010001000;
rgb[8457] = 24'b100110011001100110011001;
rgb[8458] = 24'b101010101010101010101010;
rgb[8459] = 24'b101110111011101110111011;
rgb[8460] = 24'b110011001100110011001100;
rgb[8461] = 24'b110111011101110111011101;
rgb[8462] = 24'b111011101110111011101110;
rgb[8463] = 24'b111111111111111111111111;
rgb[8464] = 24'b000000000000000000000000;
rgb[8465] = 24'b000011110001000100010010;
rgb[8466] = 24'b000111110010001100100100;
rgb[8467] = 24'b001011110011010100110110;
rgb[8468] = 24'b001111110100011101001000;
rgb[8469] = 24'b010011110101100101011010;
rgb[8470] = 24'b010111110110101001101100;
rgb[8471] = 24'b011011110111110001111110;
rgb[8472] = 24'b100000001000110110001111;
rgb[8473] = 24'b100100101001110110011111;
rgb[8474] = 24'b101001001010111010101111;
rgb[8475] = 24'b101101101011111010111111;
rgb[8476] = 24'b110010001100111011001111;
rgb[8477] = 24'b110110101101111011011111;
rgb[8478] = 24'b111011001110111011101111;
rgb[8479] = 24'b111111111111111111111111;
rgb[8480] = 24'b000000000000000000000000;
rgb[8481] = 24'b000011100001001000010011;
rgb[8482] = 24'b000111010010010100100110;
rgb[8483] = 24'b001011000011011100111001;
rgb[8484] = 24'b001110100100101001001101;
rgb[8485] = 24'b010010010101110101100000;
rgb[8486] = 24'b010110000110111101110011;
rgb[8487] = 24'b011001111000001010000110;
rgb[8488] = 24'b011110001001001110010111;
rgb[8489] = 24'b100010111010001010100110;
rgb[8490] = 24'b100111101011001010110101;
rgb[8491] = 24'b101100011100000111000100;
rgb[8492] = 24'b110001011101000011010010;
rgb[8493] = 24'b110110001110000011100001;
rgb[8494] = 24'b111010111110111111110000;
rgb[8495] = 24'b111111111111111111111111;
rgb[8496] = 24'b000000000000000000000000;
rgb[8497] = 24'b000011010001001100010100;
rgb[8498] = 24'b000110110010011000101000;
rgb[8499] = 24'b001010000011101000111101;
rgb[8500] = 24'b001101100100110101010001;
rgb[8501] = 24'b010001000110000101100101;
rgb[8502] = 24'b010100010111010001111010;
rgb[8503] = 24'b010111111000011110001110;
rgb[8504] = 24'b011100001001100110011111;
rgb[8505] = 24'b100001001010011110101101;
rgb[8506] = 24'b100110001011011010111011;
rgb[8507] = 24'b101011011100010011001000;
rgb[8508] = 24'b110000011101001111010110;
rgb[8509] = 24'b110101101110000111100011;
rgb[8510] = 24'b111010101111000011110001;
rgb[8511] = 24'b111111111111111111111111;
rgb[8512] = 24'b000000000000000000000000;
rgb[8513] = 24'b000011000001010000010101;
rgb[8514] = 24'b000110000010100000101011;
rgb[8515] = 24'b001001010011110001000000;
rgb[8516] = 24'b001100010101000001010110;
rgb[8517] = 24'b001111100110010101101011;
rgb[8518] = 24'b010010100111100110000001;
rgb[8519] = 24'b010101111000110110010110;
rgb[8520] = 24'b011010001001111010100111;
rgb[8521] = 24'b011111011010110010110100;
rgb[8522] = 24'b100100111011101011000000;
rgb[8523] = 24'b101010001100011111001101;
rgb[8524] = 24'b101111101101010111011001;
rgb[8525] = 24'b110100111110001111100110;
rgb[8526] = 24'b111010011111000111110010;
rgb[8527] = 24'b111111111111111111111111;
rgb[8528] = 24'b000000000000000000000000;
rgb[8529] = 24'b000010110001010100010110;
rgb[8530] = 24'b000101100010101000101101;
rgb[8531] = 24'b001000100011111101000100;
rgb[8532] = 24'b001011010101010001011010;
rgb[8533] = 24'b001110000110100101110001;
rgb[8534] = 24'b010001000111111010001000;
rgb[8535] = 24'b010011111001001110011110;
rgb[8536] = 24'b011000001010010010101111;
rgb[8537] = 24'b011101101011000110111011;
rgb[8538] = 24'b100011011011111011000110;
rgb[8539] = 24'b101001001100101111010001;
rgb[8540] = 24'b101110111101100011011101;
rgb[8541] = 24'b110100011110010111101000;
rgb[8542] = 24'b111010001111001011110011;
rgb[8543] = 24'b111111111111111111111111;
rgb[8544] = 24'b000000000000000000000000;
rgb[8545] = 24'b000010100001010100010111;
rgb[8546] = 24'b000101000010101100101111;
rgb[8547] = 24'b000111100100000101000111;
rgb[8548] = 24'b001010000101011101011111;
rgb[8549] = 24'b001100110110110101110110;
rgb[8550] = 24'b001111011000001110001110;
rgb[8551] = 24'b010001111001100010100110;
rgb[8552] = 24'b010110001010100110110111;
rgb[8553] = 24'b011100001011011011000001;
rgb[8554] = 24'b100001111100001011001100;
rgb[8555] = 24'b100111111100111011010110;
rgb[8556] = 24'b101101111101101011100000;
rgb[8557] = 24'b110011111110011011101010;
rgb[8558] = 24'b111001111111001011110100;
rgb[8559] = 24'b111111111111111011111110;
rgb[8560] = 24'b000000000000000000000000;
rgb[8561] = 24'b000010010001011000011000;
rgb[8562] = 24'b000100100010110100110001;
rgb[8563] = 24'b000110110100001101001010;
rgb[8564] = 24'b001001000101101001100011;
rgb[8565] = 24'b001011010111000101111100;
rgb[8566] = 24'b001101101000011110010101;
rgb[8567] = 24'b001111111001111010101110;
rgb[8568] = 24'b010100001010111110111111;
rgb[8569] = 24'b011010011011101011001000;
rgb[8570] = 24'b100000101100011011010001;
rgb[8571] = 24'b100110111101000111011010;
rgb[8572] = 24'b101101001101110011100011;
rgb[8573] = 24'b110011011110100011101100;
rgb[8574] = 24'b111001101111001111110101;
rgb[8575] = 24'b111111111111111111111111;
rgb[8576] = 24'b000000000000000000000000;
rgb[8577] = 24'b000001110001011100011010;
rgb[8578] = 24'b000011110010111000110100;
rgb[8579] = 24'b000101110100011001001110;
rgb[8580] = 24'b000111110101110101101000;
rgb[8581] = 24'b001001110111010110000010;
rgb[8582] = 24'b001011111000110010011100;
rgb[8583] = 24'b001101111010010010110110;
rgb[8584] = 24'b010010001011010111000111;
rgb[8585] = 24'b011000101011111111001111;
rgb[8586] = 24'b011111001100101011010111;
rgb[8587] = 24'b100101101101010011011111;
rgb[8588] = 24'b101100001101111111100111;
rgb[8589] = 24'b110010101110100111101111;
rgb[8590] = 24'b111001001111010011110111;
rgb[8591] = 24'b111111111111111011111110;
rgb[8592] = 24'b000000000000000000000000;
rgb[8593] = 24'b000001100001100000011011;
rgb[8594] = 24'b000011010011000000110110;
rgb[8595] = 24'b000101000100100001010001;
rgb[8596] = 24'b000110110110000101101100;
rgb[8597] = 24'b001000010111100110001000;
rgb[8598] = 24'b001010001001000110100011;
rgb[8599] = 24'b001011111010100110111110;
rgb[8600] = 24'b010000001011101011001111;
rgb[8601] = 24'b010110111100010011010110;
rgb[8602] = 24'b011101101100111011011101;
rgb[8603] = 24'b100100101101100011100011;
rgb[8604] = 24'b101011011110000111101010;
rgb[8605] = 24'b110010001110101111110001;
rgb[8606] = 24'b111000111111010111111000;
rgb[8607] = 24'b111111111111111111111111;
rgb[8608] = 24'b000000000000000000000000;
rgb[8609] = 24'b000001010001100100011100;
rgb[8610] = 24'b000010110011001000111000;
rgb[8611] = 24'b000100010100101101010101;
rgb[8612] = 24'b000101100110010001110001;
rgb[8613] = 24'b000111000111110110001101;
rgb[8614] = 24'b001000101001011010101010;
rgb[8615] = 24'b001001111010111111000110;
rgb[8616] = 24'b001110001100000011010111;
rgb[8617] = 24'b010101001100100111011101;
rgb[8618] = 24'b011100011101001011100010;
rgb[8619] = 24'b100011011101101111101000;
rgb[8620] = 24'b101010101110010011101110;
rgb[8621] = 24'b110001101110110111110011;
rgb[8622] = 24'b111000101111011011111001;
rgb[8623] = 24'b111111111111111011111110;
rgb[8624] = 24'b000000000000000000000000;
rgb[8625] = 24'b000001000001100100011101;
rgb[8626] = 24'b000010010011001100111010;
rgb[8627] = 24'b000011010100110101011000;
rgb[8628] = 24'b000100100110011101110101;
rgb[8629] = 24'b000101101000000110010011;
rgb[8630] = 24'b000110111001101110110000;
rgb[8631] = 24'b000111111011010111001110;
rgb[8632] = 24'b001100001100011011011111;
rgb[8633] = 24'b010011101100111011100011;
rgb[8634] = 24'b011010111101011011101000;
rgb[8635] = 24'b100010011101111011101100;
rgb[8636] = 24'b101001101110011011110001;
rgb[8637] = 24'b110001001110111011110101;
rgb[8638] = 24'b111000011111011011111010;
rgb[8639] = 24'b111111111111111111111111;
rgb[8640] = 24'b000000000000000000000000;
rgb[8641] = 24'b000000110001101000011110;
rgb[8642] = 24'b000001100011010100111101;
rgb[8643] = 24'b000010100101000001011011;
rgb[8644] = 24'b000011010110101001111010;
rgb[8645] = 24'b000100001000010110011001;
rgb[8646] = 24'b000101001010000010110111;
rgb[8647] = 24'b000101111011101011010110;
rgb[8648] = 24'b001010001100101111100111;
rgb[8649] = 24'b010001111101001111101010;
rgb[8650] = 24'b011001011101101011101110;
rgb[8651] = 24'b100001001110000111110001;
rgb[8652] = 24'b101000111110100111110100;
rgb[8653] = 24'b110000011111000011111000;
rgb[8654] = 24'b111000001111011111111011;
rgb[8655] = 24'b111111111111111111111111;
rgb[8656] = 24'b000000000000000000000000;
rgb[8657] = 24'b000000100001101100011111;
rgb[8658] = 24'b000001000011011100111111;
rgb[8659] = 24'b000001100101001001011111;
rgb[8660] = 24'b000010010110111001111110;
rgb[8661] = 24'b000010111000100110011110;
rgb[8662] = 24'b000011011010010110111110;
rgb[8663] = 24'b000011111100000011011110;
rgb[8664] = 24'b001000001101000111101111;
rgb[8665] = 24'b010000001101100011110001;
rgb[8666] = 24'b011000001101111011110011;
rgb[8667] = 24'b100000001110010111110101;
rgb[8668] = 24'b100111111110101111111000;
rgb[8669] = 24'b101111111111001011111010;
rgb[8670] = 24'b110111111111100011111100;
rgb[8671] = 24'b111111111111111111111111;
rgb[8672] = 24'b000000000000000000000000;
rgb[8673] = 24'b000000010001110000100000;
rgb[8674] = 24'b000000100011100001000001;
rgb[8675] = 24'b000000110101010001100010;
rgb[8676] = 24'b000001000111000110000011;
rgb[8677] = 24'b000001011000110110100100;
rgb[8678] = 24'b000001101010100111000101;
rgb[8679] = 24'b000001111100011011100110;
rgb[8680] = 24'b000110001101011111110111;
rgb[8681] = 24'b001110011101110011111000;
rgb[8682] = 24'b010110101110001011111001;
rgb[8683] = 24'b011110111110100011111010;
rgb[8684] = 24'b100111001110110111111011;
rgb[8685] = 24'b101111011111001111111100;
rgb[8686] = 24'b110111101111100111111101;
rgb[8687] = 24'b111111111111111111111111;
rgb[8688] = 24'b000000000000000000000000;
rgb[8689] = 24'b000000000001110100100010;
rgb[8690] = 24'b000000000011101001000100;
rgb[8691] = 24'b000000000101011101100110;
rgb[8692] = 24'b000000000111010010001000;
rgb[8693] = 24'b000000001001000110101010;
rgb[8694] = 24'b000000001010111011001100;
rgb[8695] = 24'b000000001100101111101110;
rgb[8696] = 24'b000100011101110011111110;
rgb[8697] = 24'b001100101110000111111111;
rgb[8698] = 24'b010101011110011011111110;
rgb[8699] = 24'b011101101110101111111111;
rgb[8700] = 24'b100110011111000011111111;
rgb[8701] = 24'b101110111111010111111111;
rgb[8702] = 24'b110111011111101011111111;
rgb[8703] = 24'b111111111111111111111111;
rgb[8704] = 24'b000000000000000000000000;
rgb[8705] = 24'b000100010001000100010001;
rgb[8706] = 24'b001000100010001000100010;
rgb[8707] = 24'b001100110011001100110011;
rgb[8708] = 24'b010001000100010001000100;
rgb[8709] = 24'b010101010101010101010101;
rgb[8710] = 24'b011001100110011001100110;
rgb[8711] = 24'b011101110111011101110111;
rgb[8712] = 24'b100010001000100010001000;
rgb[8713] = 24'b100110011001100110011001;
rgb[8714] = 24'b101010101010101010101010;
rgb[8715] = 24'b101110111011101110111011;
rgb[8716] = 24'b110011001100110011001100;
rgb[8717] = 24'b110111011101110111011101;
rgb[8718] = 24'b111011101110111011101110;
rgb[8719] = 24'b111111111111111111111111;
rgb[8720] = 24'b000000000000000000000000;
rgb[8721] = 24'b000011110001000100010010;
rgb[8722] = 24'b000111110010001100100100;
rgb[8723] = 24'b001011110011010000110110;
rgb[8724] = 24'b001111110100011001001000;
rgb[8725] = 24'b010011110101011101011010;
rgb[8726] = 24'b010111110110100101101100;
rgb[8727] = 24'b011011110111101101111110;
rgb[8728] = 24'b100000001000110010001111;
rgb[8729] = 24'b100100101001110010011111;
rgb[8730] = 24'b101001001010110010101111;
rgb[8731] = 24'b101101101011110110111111;
rgb[8732] = 24'b110010001100110111001111;
rgb[8733] = 24'b110110101101111011011111;
rgb[8734] = 24'b111011001110111011101111;
rgb[8735] = 24'b111111111111111111111111;
rgb[8736] = 24'b000000000000000000000000;
rgb[8737] = 24'b000011100001001000010011;
rgb[8738] = 24'b000111010010010000100110;
rgb[8739] = 24'b001011000011011000111001;
rgb[8740] = 24'b001110100100100001001101;
rgb[8741] = 24'b010010010101101001100000;
rgb[8742] = 24'b010110000110110101110011;
rgb[8743] = 24'b011001110111111110000110;
rgb[8744] = 24'b011110001001000010010111;
rgb[8745] = 24'b100010111010000010100110;
rgb[8746] = 24'b100111101010111110110101;
rgb[8747] = 24'b101100011011111111000100;
rgb[8748] = 24'b110001011100111111010010;
rgb[8749] = 24'b110110001101111111100001;
rgb[8750] = 24'b111010111110111111110000;
rgb[8751] = 24'b111111111111111111111111;
rgb[8752] = 24'b000000000000000000000000;
rgb[8753] = 24'b000011010001001000010100;
rgb[8754] = 24'b000110110010010100101000;
rgb[8755] = 24'b001010000011100000111101;
rgb[8756] = 24'b001101100100101101010001;
rgb[8757] = 24'b010001000101110101100101;
rgb[8758] = 24'b010100010111000001111010;
rgb[8759] = 24'b010111111000001110001110;
rgb[8760] = 24'b011100001001010010011111;
rgb[8761] = 24'b100001001010001110101101;
rgb[8762] = 24'b100110001011001010111011;
rgb[8763] = 24'b101011011100001011001000;
rgb[8764] = 24'b110000011101000111010110;
rgb[8765] = 24'b110101101110000011100011;
rgb[8766] = 24'b111010101110111111110001;
rgb[8767] = 24'b111111111111111111111111;
rgb[8768] = 24'b000000000000000000000000;
rgb[8769] = 24'b000011000001001100010101;
rgb[8770] = 24'b000110000010011000101011;
rgb[8771] = 24'b001001010011101001000000;
rgb[8772] = 24'b001100010100110101010110;
rgb[8773] = 24'b001111100110000001101011;
rgb[8774] = 24'b010010100111010010000001;
rgb[8775] = 24'b010101111000011110010110;
rgb[8776] = 24'b011010001001100010100111;
rgb[8777] = 24'b011111011010011110110100;
rgb[8778] = 24'b100100111011010111000000;
rgb[8779] = 24'b101010001100010011001101;
rgb[8780] = 24'b101111101101001111011001;
rgb[8781] = 24'b110100111110000111100110;
rgb[8782] = 24'b111010011111000011110010;
rgb[8783] = 24'b111111111111111111111111;
rgb[8784] = 24'b000000000000000000000000;
rgb[8785] = 24'b000010110001001100010110;
rgb[8786] = 24'b000101100010011100101101;
rgb[8787] = 24'b001000100011101101000100;
rgb[8788] = 24'b001011010100111101011010;
rgb[8789] = 24'b001110000110001101110001;
rgb[8790] = 24'b010001000111011110001000;
rgb[8791] = 24'b010011111000101110011110;
rgb[8792] = 24'b011000001001110010101111;
rgb[8793] = 24'b011101101010101010111011;
rgb[8794] = 24'b100011011011100011000110;
rgb[8795] = 24'b101001001100011011010001;
rgb[8796] = 24'b101110111101010011011101;
rgb[8797] = 24'b110100011110001011101000;
rgb[8798] = 24'b111010001111000011110011;
rgb[8799] = 24'b111111111111111111111111;
rgb[8800] = 24'b000000000000000000000000;
rgb[8801] = 24'b000010100001010000010111;
rgb[8802] = 24'b000101000010100100101111;
rgb[8803] = 24'b000111100011110101000111;
rgb[8804] = 24'b001010000101001001011111;
rgb[8805] = 24'b001100110110011001110110;
rgb[8806] = 24'b001111010111101110001110;
rgb[8807] = 24'b010001111000111110100110;
rgb[8808] = 24'b010110001010000010110111;
rgb[8809] = 24'b011100001010111011000001;
rgb[8810] = 24'b100001111011101111001100;
rgb[8811] = 24'b100111111100100111010110;
rgb[8812] = 24'b101101111101011011100000;
rgb[8813] = 24'b110011111110010011101010;
rgb[8814] = 24'b111001111111000111110100;
rgb[8815] = 24'b111111111111111011111110;
rgb[8816] = 24'b000000000000000000000000;
rgb[8817] = 24'b000010010001010100011000;
rgb[8818] = 24'b000100100010101000110001;
rgb[8819] = 24'b000110110011111101001010;
rgb[8820] = 24'b001001000101010001100011;
rgb[8821] = 24'b001011010110100101111100;
rgb[8822] = 24'b001101100111111010010101;
rgb[8823] = 24'b001111111001010010101110;
rgb[8824] = 24'b010100001010010110111111;
rgb[8825] = 24'b011010011011000111001000;
rgb[8826] = 24'b100000101011111011010001;
rgb[8827] = 24'b100110111100101111011010;
rgb[8828] = 24'b101101001101100011100011;
rgb[8829] = 24'b110011011110010111101100;
rgb[8830] = 24'b111001101111001011110101;
rgb[8831] = 24'b111111111111111111111111;
rgb[8832] = 24'b000000000000000000000000;
rgb[8833] = 24'b000001110001010100011010;
rgb[8834] = 24'b000011110010101100110100;
rgb[8835] = 24'b000101110100000101001110;
rgb[8836] = 24'b000111110101011001101000;
rgb[8837] = 24'b001001110110110010000010;
rgb[8838] = 24'b001011111000001010011100;
rgb[8839] = 24'b001101111001100010110110;
rgb[8840] = 24'b010010001010100111000111;
rgb[8841] = 24'b011000101011010111001111;
rgb[8842] = 24'b011111001100000111010111;
rgb[8843] = 24'b100101101100110111011111;
rgb[8844] = 24'b101100001101101011100111;
rgb[8845] = 24'b110010101110011011101111;
rgb[8846] = 24'b111001001111001011110111;
rgb[8847] = 24'b111111111111111011111110;
rgb[8848] = 24'b000000000000000000000000;
rgb[8849] = 24'b000001100001011000011011;
rgb[8850] = 24'b000011010010110000110110;
rgb[8851] = 24'b000101000100001101010001;
rgb[8852] = 24'b000110110101100101101100;
rgb[8853] = 24'b001000010110111110001000;
rgb[8854] = 24'b001010001000011010100011;
rgb[8855] = 24'b001011111001110010111110;
rgb[8856] = 24'b010000001010110111001111;
rgb[8857] = 24'b010110111011100111010110;
rgb[8858] = 24'b011101101100010011011101;
rgb[8859] = 24'b100100101101000011100011;
rgb[8860] = 24'b101011011101110011101010;
rgb[8861] = 24'b110010001110011111110001;
rgb[8862] = 24'b111000111111001111111000;
rgb[8863] = 24'b111111111111111111111111;
rgb[8864] = 24'b000000000000000000000000;
rgb[8865] = 24'b000001010001011000011100;
rgb[8866] = 24'b000010110010110100111000;
rgb[8867] = 24'b000100010100010001010101;
rgb[8868] = 24'b000101100101101101110001;
rgb[8869] = 24'b000111000111001010001101;
rgb[8870] = 24'b001000101000100110101010;
rgb[8871] = 24'b001001111010000011000110;
rgb[8872] = 24'b001110001011000111010111;
rgb[8873] = 24'b010101001011110011011101;
rgb[8874] = 24'b011100011100011111100010;
rgb[8875] = 24'b100011011101001011101000;
rgb[8876] = 24'b101010101101110111101110;
rgb[8877] = 24'b110001101110100011110011;
rgb[8878] = 24'b111000101111001111111001;
rgb[8879] = 24'b111111111111111011111110;
rgb[8880] = 24'b000000000000000000000000;
rgb[8881] = 24'b000001000001011100011101;
rgb[8882] = 24'b000010010010111100111010;
rgb[8883] = 24'b000011010100011001011000;
rgb[8884] = 24'b000100100101111001110101;
rgb[8885] = 24'b000101100111010110010011;
rgb[8886] = 24'b000110111000110110110000;
rgb[8887] = 24'b000111111010010011001110;
rgb[8888] = 24'b001100001011010111011111;
rgb[8889] = 24'b010011101100000011100011;
rgb[8890] = 24'b011010111100101011101000;
rgb[8891] = 24'b100010011101010111101100;
rgb[8892] = 24'b101001101101111111110001;
rgb[8893] = 24'b110001001110101011110101;
rgb[8894] = 24'b111000011111010011111010;
rgb[8895] = 24'b111111111111111111111111;
rgb[8896] = 24'b000000000000000000000000;
rgb[8897] = 24'b000000110001100000011110;
rgb[8898] = 24'b000001100011000000111101;
rgb[8899] = 24'b000010100100100001011011;
rgb[8900] = 24'b000011010110000001111010;
rgb[8901] = 24'b000100000111100010011001;
rgb[8902] = 24'b000101001001000010110111;
rgb[8903] = 24'b000101111010100011010110;
rgb[8904] = 24'b001010001011100111100111;
rgb[8905] = 24'b010001111100001111101010;
rgb[8906] = 24'b011001011100110111101110;
rgb[8907] = 24'b100001001101011111110001;
rgb[8908] = 24'b101000111110000111110100;
rgb[8909] = 24'b110000011110101111111000;
rgb[8910] = 24'b111000001111010111111011;
rgb[8911] = 24'b111111111111111111111111;
rgb[8912] = 24'b000000000000000000000000;
rgb[8913] = 24'b000000100001100000011111;
rgb[8914] = 24'b000001000011000100111111;
rgb[8915] = 24'b000001100100101001011111;
rgb[8916] = 24'b000010010110001001111110;
rgb[8917] = 24'b000010110111101110011110;
rgb[8918] = 24'b000011011001010010111110;
rgb[8919] = 24'b000011111010110111011110;
rgb[8920] = 24'b001000001011111011101111;
rgb[8921] = 24'b010000001100011111110001;
rgb[8922] = 24'b011000001101000011110011;
rgb[8923] = 24'b100000001101100111110101;
rgb[8924] = 24'b100111111110001111111000;
rgb[8925] = 24'b101111111110110011111010;
rgb[8926] = 24'b110111111111010111111100;
rgb[8927] = 24'b111111111111111111111111;
rgb[8928] = 24'b000000000000000000000000;
rgb[8929] = 24'b000000010001100100100000;
rgb[8930] = 24'b000000100011001001000001;
rgb[8931] = 24'b000000110100101101100010;
rgb[8932] = 24'b000001000110010110000011;
rgb[8933] = 24'b000001010111111010100100;
rgb[8934] = 24'b000001101001011111000101;
rgb[8935] = 24'b000001111011000111100110;
rgb[8936] = 24'b000110001100001011110111;
rgb[8937] = 24'b001110011100101011111000;
rgb[8938] = 24'b010110101101001111111001;
rgb[8939] = 24'b011110111101110011111010;
rgb[8940] = 24'b100111001110010011111011;
rgb[8941] = 24'b101111011110110111111100;
rgb[8942] = 24'b110111101111011011111101;
rgb[8943] = 24'b111111111111111111111111;
rgb[8944] = 24'b000000000000000000000000;
rgb[8945] = 24'b000000000001100100100010;
rgb[8946] = 24'b000000000011001101000100;
rgb[8947] = 24'b000000000100110101100110;
rgb[8948] = 24'b000000000110011110001000;
rgb[8949] = 24'b000000001000000110101010;
rgb[8950] = 24'b000000001001101111001100;
rgb[8951] = 24'b000000001011010111101110;
rgb[8952] = 24'b000100011100011011111110;
rgb[8953] = 24'b001100101100111011111111;
rgb[8954] = 24'b010101011101011011111110;
rgb[8955] = 24'b011101101101111011111111;
rgb[8956] = 24'b100110011110011011111111;
rgb[8957] = 24'b101110111110111011111111;
rgb[8958] = 24'b110111011111011011111111;
rgb[8959] = 24'b111111111111111111111111;
rgb[8960] = 24'b000000000000000000000000;
rgb[8961] = 24'b000100010001000100010001;
rgb[8962] = 24'b001000100010001000100010;
rgb[8963] = 24'b001100110011001100110011;
rgb[8964] = 24'b010001000100010001000100;
rgb[8965] = 24'b010101010101010101010101;
rgb[8966] = 24'b011001100110011001100110;
rgb[8967] = 24'b011101110111011101110111;
rgb[8968] = 24'b100010001000100010001000;
rgb[8969] = 24'b100110011001100110011001;
rgb[8970] = 24'b101010101010101010101010;
rgb[8971] = 24'b101110111011101110111011;
rgb[8972] = 24'b110011001100110011001100;
rgb[8973] = 24'b110111011101110111011101;
rgb[8974] = 24'b111011101110111011101110;
rgb[8975] = 24'b111111111111111111111111;
rgb[8976] = 24'b000000000000000000000000;
rgb[8977] = 24'b000011110001000100010010;
rgb[8978] = 24'b000111110010001000100100;
rgb[8979] = 24'b001011110011010000110110;
rgb[8980] = 24'b001111110100010101001000;
rgb[8981] = 24'b010011110101011001011010;
rgb[8982] = 24'b010111110110100001101100;
rgb[8983] = 24'b011011110111100101111110;
rgb[8984] = 24'b100000001000101010001111;
rgb[8985] = 24'b100100101001101110011111;
rgb[8986] = 24'b101001001010101110101111;
rgb[8987] = 24'b101101101011110010111111;
rgb[8988] = 24'b110010001100110111001111;
rgb[8989] = 24'b110110101101110111011111;
rgb[8990] = 24'b111011001110111011101111;
rgb[8991] = 24'b111111111111111111111111;
rgb[8992] = 24'b000000000000000000000000;
rgb[8993] = 24'b000011100001000100010011;
rgb[8994] = 24'b000111010010001100100110;
rgb[8995] = 24'b001011000011010100111001;
rgb[8996] = 24'b001110100100011101001101;
rgb[8997] = 24'b010010010101100001100000;
rgb[8998] = 24'b010110000110101001110011;
rgb[8999] = 24'b011001110111110010000110;
rgb[9000] = 24'b011110001000110110010111;
rgb[9001] = 24'b100010111001110110100110;
rgb[9002] = 24'b100111101010110110110101;
rgb[9003] = 24'b101100011011111011000100;
rgb[9004] = 24'b110001011100111011010010;
rgb[9005] = 24'b110110001101111011100001;
rgb[9006] = 24'b111010111110111011110000;
rgb[9007] = 24'b111111111111111111111111;
rgb[9008] = 24'b000000000000000000000000;
rgb[9009] = 24'b000011010001001000010100;
rgb[9010] = 24'b000110110010010000101000;
rgb[9011] = 24'b001010000011011000111101;
rgb[9012] = 24'b001101100100100001010001;
rgb[9013] = 24'b010001000101101001100101;
rgb[9014] = 24'b010100010110110001111010;
rgb[9015] = 24'b010111110111111010001110;
rgb[9016] = 24'b011100001000111110011111;
rgb[9017] = 24'b100001001001111110101101;
rgb[9018] = 24'b100110001010111110111011;
rgb[9019] = 24'b101011011011111111001000;
rgb[9020] = 24'b110000011100111111010110;
rgb[9021] = 24'b110101101101111111100011;
rgb[9022] = 24'b111010101110111111110001;
rgb[9023] = 24'b111111111111111111111111;
rgb[9024] = 24'b000000000000000000000000;
rgb[9025] = 24'b000011000001001000010101;
rgb[9026] = 24'b000110000010010100101011;
rgb[9027] = 24'b001001010011011101000000;
rgb[9028] = 24'b001100010100101001010110;
rgb[9029] = 24'b001111100101110001101011;
rgb[9030] = 24'b010010100110111110000001;
rgb[9031] = 24'b010101111000000110010110;
rgb[9032] = 24'b011010001001001010100111;
rgb[9033] = 24'b011111011010001010110100;
rgb[9034] = 24'b100100111011000111000000;
rgb[9035] = 24'b101010001100000111001101;
rgb[9036] = 24'b101111101101000011011001;
rgb[9037] = 24'b110100111110000011100110;
rgb[9038] = 24'b111010011110111111110010;
rgb[9039] = 24'b111111111111111111111111;
rgb[9040] = 24'b000000000000000000000000;
rgb[9041] = 24'b000010110001001000010110;
rgb[9042] = 24'b000101100010010100101101;
rgb[9043] = 24'b001000100011100001000100;
rgb[9044] = 24'b001011010100101101011010;
rgb[9045] = 24'b001110000101111001110001;
rgb[9046] = 24'b010001000111000110001000;
rgb[9047] = 24'b010011111000010010011110;
rgb[9048] = 24'b011000001001010110101111;
rgb[9049] = 24'b011101101010010010111011;
rgb[9050] = 24'b100011011011001111000110;
rgb[9051] = 24'b101001001100001011010001;
rgb[9052] = 24'b101110111101000111011101;
rgb[9053] = 24'b110100011110000011101000;
rgb[9054] = 24'b111010001110111111110011;
rgb[9055] = 24'b111111111111111111111111;
rgb[9056] = 24'b000000000000000000000000;
rgb[9057] = 24'b000010100001001100010111;
rgb[9058] = 24'b000101000010011000101111;
rgb[9059] = 24'b000111100011100101000111;
rgb[9060] = 24'b001010000100110101011111;
rgb[9061] = 24'b001100110110000001110110;
rgb[9062] = 24'b001111010111001110001110;
rgb[9063] = 24'b010001111000011010100110;
rgb[9064] = 24'b010110001001011110110111;
rgb[9065] = 24'b011100001010011011000001;
rgb[9066] = 24'b100001111011010111001100;
rgb[9067] = 24'b100111111100010011010110;
rgb[9068] = 24'b101101111101001011100000;
rgb[9069] = 24'b110011111110000111101010;
rgb[9070] = 24'b111001111111000011110100;
rgb[9071] = 24'b111111111111111011111110;
rgb[9072] = 24'b000000000000000000000000;
rgb[9073] = 24'b000010010001001100011000;
rgb[9074] = 24'b000100100010011100110001;
rgb[9075] = 24'b000110110011101001001010;
rgb[9076] = 24'b001001000100111001100011;
rgb[9077] = 24'b001011010110001001111100;
rgb[9078] = 24'b001101100111010110010101;
rgb[9079] = 24'b001111111000100110101110;
rgb[9080] = 24'b010100001001101010111111;
rgb[9081] = 24'b011010011010100011001000;
rgb[9082] = 24'b100000101011011111010001;
rgb[9083] = 24'b100110111100010111011010;
rgb[9084] = 24'b101101001101001111100011;
rgb[9085] = 24'b110011011110001011101100;
rgb[9086] = 24'b111001101111000011110101;
rgb[9087] = 24'b111111111111111111111111;
rgb[9088] = 24'b000000000000000000000000;
rgb[9089] = 24'b000001110001010000011010;
rgb[9090] = 24'b000011110010100000110100;
rgb[9091] = 24'b000101110011110001001110;
rgb[9092] = 24'b000111110101000001101000;
rgb[9093] = 24'b001001110110010010000010;
rgb[9094] = 24'b001011110111100010011100;
rgb[9095] = 24'b001101111000110010110110;
rgb[9096] = 24'b010010001001110111000111;
rgb[9097] = 24'b011000101010101111001111;
rgb[9098] = 24'b011111001011100111010111;
rgb[9099] = 24'b100101101100011111011111;
rgb[9100] = 24'b101100001101010111100111;
rgb[9101] = 24'b110010101110001111101111;
rgb[9102] = 24'b111001001111000111110111;
rgb[9103] = 24'b111111111111111011111110;
rgb[9104] = 24'b000000000000000000000000;
rgb[9105] = 24'b000001100001010000011011;
rgb[9106] = 24'b000011010010100000110110;
rgb[9107] = 24'b000101000011110101010001;
rgb[9108] = 24'b000110110101000101101100;
rgb[9109] = 24'b001000010110010110001000;
rgb[9110] = 24'b001010000111101010100011;
rgb[9111] = 24'b001011111000111010111110;
rgb[9112] = 24'b010000001001111111001111;
rgb[9113] = 24'b010110111010110111010110;
rgb[9114] = 24'b011101101011101011011101;
rgb[9115] = 24'b100100101100100011100011;
rgb[9116] = 24'b101011011101011011101010;
rgb[9117] = 24'b110010001110001111110001;
rgb[9118] = 24'b111000111111000111111000;
rgb[9119] = 24'b111111111111111111111111;
rgb[9120] = 24'b000000000000000000000000;
rgb[9121] = 24'b000001010001010000011100;
rgb[9122] = 24'b000010110010100100111000;
rgb[9123] = 24'b000100010011111001010101;
rgb[9124] = 24'b000101100101001101110001;
rgb[9125] = 24'b000111000110011110001101;
rgb[9126] = 24'b001000100111110010101010;
rgb[9127] = 24'b001001111001000111000110;
rgb[9128] = 24'b001110001010001011010111;
rgb[9129] = 24'b010101001010111111011101;
rgb[9130] = 24'b011100011011110011100010;
rgb[9131] = 24'b100011011100101011101000;
rgb[9132] = 24'b101010101101011111101110;
rgb[9133] = 24'b110001101110010011110011;
rgb[9134] = 24'b111000101111000111111001;
rgb[9135] = 24'b111111111111111011111110;
rgb[9136] = 24'b000000000000000000000000;
rgb[9137] = 24'b000001000001010100011101;
rgb[9138] = 24'b000010010010101000111010;
rgb[9139] = 24'b000011010011111101011000;
rgb[9140] = 24'b000100100101010001110101;
rgb[9141] = 24'b000101100110100110010011;
rgb[9142] = 24'b000110110111111010110000;
rgb[9143] = 24'b000111111001010011001110;
rgb[9144] = 24'b001100001010010111011111;
rgb[9145] = 24'b010011101011000111100011;
rgb[9146] = 24'b011010111011111011101000;
rgb[9147] = 24'b100010011100101111101100;
rgb[9148] = 24'b101001101101100011110001;
rgb[9149] = 24'b110001001110010111110101;
rgb[9150] = 24'b111000011111001011111010;
rgb[9151] = 24'b111111111111111111111111;
rgb[9152] = 24'b000000000000000000000000;
rgb[9153] = 24'b000000110001010100011110;
rgb[9154] = 24'b000001100010101100111101;
rgb[9155] = 24'b000010100100000001011011;
rgb[9156] = 24'b000011010101011001111010;
rgb[9157] = 24'b000100000110101110011001;
rgb[9158] = 24'b000101001000000110110111;
rgb[9159] = 24'b000101111001011011010110;
rgb[9160] = 24'b001010001010011111100111;
rgb[9161] = 24'b010001111011010011101010;
rgb[9162] = 24'b011001011100000011101110;
rgb[9163] = 24'b100001001100110111110001;
rgb[9164] = 24'b101000111101100111110100;
rgb[9165] = 24'b110000011110011011111000;
rgb[9166] = 24'b111000001111001011111011;
rgb[9167] = 24'b111111111111111111111111;
rgb[9168] = 24'b000000000000000000000000;
rgb[9169] = 24'b000000100001010100011111;
rgb[9170] = 24'b000001000010101100111111;
rgb[9171] = 24'b000001100100000101011111;
rgb[9172] = 24'b000010010101011101111110;
rgb[9173] = 24'b000010110110110110011110;
rgb[9174] = 24'b000011011000001110111110;
rgb[9175] = 24'b000011111001100111011110;
rgb[9176] = 24'b001000001010101011101111;
rgb[9177] = 24'b010000001011011011110001;
rgb[9178] = 24'b011000001100001011110011;
rgb[9179] = 24'b100000001100111011110101;
rgb[9180] = 24'b100111111101101011111000;
rgb[9181] = 24'b101111111110011011111010;
rgb[9182] = 24'b110111111111001011111100;
rgb[9183] = 24'b111111111111111111111111;
rgb[9184] = 24'b000000000000000000000000;
rgb[9185] = 24'b000000010001011000100000;
rgb[9186] = 24'b000000100010110001000001;
rgb[9187] = 24'b000000110100001001100010;
rgb[9188] = 24'b000001000101100110000011;
rgb[9189] = 24'b000001010110111110100100;
rgb[9190] = 24'b000001101000010111000101;
rgb[9191] = 24'b000001111001110011100110;
rgb[9192] = 24'b000110001010110111110111;
rgb[9193] = 24'b001110011011100011111000;
rgb[9194] = 24'b010110101100010011111001;
rgb[9195] = 24'b011110111101000011111010;
rgb[9196] = 24'b100111001101101111111011;
rgb[9197] = 24'b101111011110011111111100;
rgb[9198] = 24'b110111101111001111111101;
rgb[9199] = 24'b111111111111111111111111;
rgb[9200] = 24'b000000000000000000000000;
rgb[9201] = 24'b000000000001011000100010;
rgb[9202] = 24'b000000000010110101000100;
rgb[9203] = 24'b000000000100001101100110;
rgb[9204] = 24'b000000000101101010001000;
rgb[9205] = 24'b000000000111000110101010;
rgb[9206] = 24'b000000001000011111001100;
rgb[9207] = 24'b000000001001111011101110;
rgb[9208] = 24'b000100011010111111111110;
rgb[9209] = 24'b001100101011101011111111;
rgb[9210] = 24'b010101011100011011111110;
rgb[9211] = 24'b011101101101000111111111;
rgb[9212] = 24'b100110011101110011111111;
rgb[9213] = 24'b101110111110100011111111;
rgb[9214] = 24'b110111011111001111111111;
rgb[9215] = 24'b111111111111111111111111;
rgb[9216] = 24'b000000000000000000000000;
rgb[9217] = 24'b000100010001000100010001;
rgb[9218] = 24'b001000100010001000100010;
rgb[9219] = 24'b001100110011001100110011;
rgb[9220] = 24'b010001000100010001000100;
rgb[9221] = 24'b010101010101010101010101;
rgb[9222] = 24'b011001100110011001100110;
rgb[9223] = 24'b011101110111011101110111;
rgb[9224] = 24'b100010001000100010001000;
rgb[9225] = 24'b100110011001100110011001;
rgb[9226] = 24'b101010101010101010101010;
rgb[9227] = 24'b101110111011101110111011;
rgb[9228] = 24'b110011001100110011001100;
rgb[9229] = 24'b110111011101110111011101;
rgb[9230] = 24'b111011101110111011101110;
rgb[9231] = 24'b111111111111111111111111;
rgb[9232] = 24'b000000000000000000000000;
rgb[9233] = 24'b000011110001000100010010;
rgb[9234] = 24'b000111110010001000100100;
rgb[9235] = 24'b001011110011001100110110;
rgb[9236] = 24'b001111110100010001001000;
rgb[9237] = 24'b010011110101010101011010;
rgb[9238] = 24'b010111110110011001101100;
rgb[9239] = 24'b011011110111100001111110;
rgb[9240] = 24'b100000001000100110001111;
rgb[9241] = 24'b100100101001100110011111;
rgb[9242] = 24'b101001001010101010101111;
rgb[9243] = 24'b101101101011101110111111;
rgb[9244] = 24'b110010001100110011001111;
rgb[9245] = 24'b110110101101110111011111;
rgb[9246] = 24'b111011001110111011101111;
rgb[9247] = 24'b111111111111111111111111;
rgb[9248] = 24'b000000000000000000000000;
rgb[9249] = 24'b000011100001000100010011;
rgb[9250] = 24'b000111010010001000100110;
rgb[9251] = 24'b001011000011001100111001;
rgb[9252] = 24'b001110100100010101001101;
rgb[9253] = 24'b010010010101011001100000;
rgb[9254] = 24'b010110000110011101110011;
rgb[9255] = 24'b011001110111100110000110;
rgb[9256] = 24'b011110001000101010010111;
rgb[9257] = 24'b100010111001101010100110;
rgb[9258] = 24'b100111101010101110110101;
rgb[9259] = 24'b101100011011110011000100;
rgb[9260] = 24'b110001011100110011010010;
rgb[9261] = 24'b110110001101110111100001;
rgb[9262] = 24'b111010111110111011110000;
rgb[9263] = 24'b111111111111111111111111;
rgb[9264] = 24'b000000000000000000000000;
rgb[9265] = 24'b000011010001000100010100;
rgb[9266] = 24'b000110110010001000101000;
rgb[9267] = 24'b001010000011010000111101;
rgb[9268] = 24'b001101100100010101010001;
rgb[9269] = 24'b010001000101011101100101;
rgb[9270] = 24'b010100010110100001111010;
rgb[9271] = 24'b010111110111101010001110;
rgb[9272] = 24'b011100001000101110011111;
rgb[9273] = 24'b100001001001101110101101;
rgb[9274] = 24'b100110001010110010111011;
rgb[9275] = 24'b101011011011110011001000;
rgb[9276] = 24'b110000011100110111010110;
rgb[9277] = 24'b110101101101110111100011;
rgb[9278] = 24'b111010101110111011110001;
rgb[9279] = 24'b111111111111111111111111;
rgb[9280] = 24'b000000000000000000000000;
rgb[9281] = 24'b000011000001000100010101;
rgb[9282] = 24'b000110000010001100101011;
rgb[9283] = 24'b001001010011010001000000;
rgb[9284] = 24'b001100010100011001010110;
rgb[9285] = 24'b001111100101100001101011;
rgb[9286] = 24'b010010100110100110000001;
rgb[9287] = 24'b010101110111101110010110;
rgb[9288] = 24'b011010001000110010100111;
rgb[9289] = 24'b011111011001110010110100;
rgb[9290] = 24'b100100111010110111000000;
rgb[9291] = 24'b101010001011110111001101;
rgb[9292] = 24'b101111101100110111011001;
rgb[9293] = 24'b110100111101111011100110;
rgb[9294] = 24'b111010011110111011110010;
rgb[9295] = 24'b111111111111111111111111;
rgb[9296] = 24'b000000000000000000000000;
rgb[9297] = 24'b000010110001000100010110;
rgb[9298] = 24'b000101100010001100101101;
rgb[9299] = 24'b001000100011010101000100;
rgb[9300] = 24'b001011010100011101011010;
rgb[9301] = 24'b001110000101100101110001;
rgb[9302] = 24'b010001000110101010001000;
rgb[9303] = 24'b010011110111110010011110;
rgb[9304] = 24'b011000001000110110101111;
rgb[9305] = 24'b011101101001110110111011;
rgb[9306] = 24'b100011011010111011000110;
rgb[9307] = 24'b101001001011111011010001;
rgb[9308] = 24'b101110111100111011011101;
rgb[9309] = 24'b110100011101111011101000;
rgb[9310] = 24'b111010001110111011110011;
rgb[9311] = 24'b111111111111111111111111;
rgb[9312] = 24'b000000000000000000000000;
rgb[9313] = 24'b000010100001000100010111;
rgb[9314] = 24'b000101000010001100101111;
rgb[9315] = 24'b000111100011010101000111;
rgb[9316] = 24'b001010000100011101011111;
rgb[9317] = 24'b001100110101100101110110;
rgb[9318] = 24'b001111010110101110001110;
rgb[9319] = 24'b010001110111110110100110;
rgb[9320] = 24'b010110001000111010110111;
rgb[9321] = 24'b011100001001111011000001;
rgb[9322] = 24'b100001111010111011001100;
rgb[9323] = 24'b100111111011111011010110;
rgb[9324] = 24'b101101111100111011100000;
rgb[9325] = 24'b110011111101111011101010;
rgb[9326] = 24'b111001111110111011110100;
rgb[9327] = 24'b111111111111111011111110;
rgb[9328] = 24'b000000000000000000000000;
rgb[9329] = 24'b000010010001001000011000;
rgb[9330] = 24'b000100100010010000110001;
rgb[9331] = 24'b000110110011011001001010;
rgb[9332] = 24'b001001000100100001100011;
rgb[9333] = 24'b001011010101101001111100;
rgb[9334] = 24'b001101100110110010010101;
rgb[9335] = 24'b001111110111111010101110;
rgb[9336] = 24'b010100001000111110111111;
rgb[9337] = 24'b011010011001111111001000;
rgb[9338] = 24'b100000101010111111010001;
rgb[9339] = 24'b100110111011111111011010;
rgb[9340] = 24'b101101001100111111100011;
rgb[9341] = 24'b110011011101111111101100;
rgb[9342] = 24'b111001101110111111110101;
rgb[9343] = 24'b111111111111111111111111;
rgb[9344] = 24'b000000000000000000000000;
rgb[9345] = 24'b000001110001001000011010;
rgb[9346] = 24'b000011110010010000110100;
rgb[9347] = 24'b000101110011011001001110;
rgb[9348] = 24'b000111110100100101101000;
rgb[9349] = 24'b001001110101101110000010;
rgb[9350] = 24'b001011110110110110011100;
rgb[9351] = 24'b001101111000000010110110;
rgb[9352] = 24'b010010001001000111000111;
rgb[9353] = 24'b011000101010000011001111;
rgb[9354] = 24'b011111001011000011010111;
rgb[9355] = 24'b100101101100000011011111;
rgb[9356] = 24'b101100001100111111100111;
rgb[9357] = 24'b110010101101111111101111;
rgb[9358] = 24'b111001001110111111110111;
rgb[9359] = 24'b111111111111111011111110;
rgb[9360] = 24'b000000000000000000000000;
rgb[9361] = 24'b000001100001001000011011;
rgb[9362] = 24'b000011010010010000110110;
rgb[9363] = 24'b000101000011011101010001;
rgb[9364] = 24'b000110110100100101101100;
rgb[9365] = 24'b001000010101110010001000;
rgb[9366] = 24'b001010000110111010100011;
rgb[9367] = 24'b001011111000000110111110;
rgb[9368] = 24'b010000001001001011001111;
rgb[9369] = 24'b010110111010000111010110;
rgb[9370] = 24'b011101101011000111011101;
rgb[9371] = 24'b100100101100000011100011;
rgb[9372] = 24'b101011011101000011101010;
rgb[9373] = 24'b110010001101111111110001;
rgb[9374] = 24'b111000111110111111111000;
rgb[9375] = 24'b111111111111111111111111;
rgb[9376] = 24'b000000000000000000000000;
rgb[9377] = 24'b000001010001001000011100;
rgb[9378] = 24'b000010110010010100111000;
rgb[9379] = 24'b000100010011011101010101;
rgb[9380] = 24'b000101100100101001110001;
rgb[9381] = 24'b000111000101110110001101;
rgb[9382] = 24'b001000100110111110101010;
rgb[9383] = 24'b001001111000001011000110;
rgb[9384] = 24'b001110001001001111010111;
rgb[9385] = 24'b010101001010001011011101;
rgb[9386] = 24'b011100011011001011100010;
rgb[9387] = 24'b100011011100000111101000;
rgb[9388] = 24'b101010101101000011101110;
rgb[9389] = 24'b110001101110000011110011;
rgb[9390] = 24'b111000101110111111111001;
rgb[9391] = 24'b111111111111111011111110;
rgb[9392] = 24'b000000000000000000000000;
rgb[9393] = 24'b000001000001001000011101;
rgb[9394] = 24'b000010010010010100111010;
rgb[9395] = 24'b000011010011100001011000;
rgb[9396] = 24'b000100100100101101110101;
rgb[9397] = 24'b000101100101110110010011;
rgb[9398] = 24'b000110110111000010110000;
rgb[9399] = 24'b000111111000001111001110;
rgb[9400] = 24'b001100001001010011011111;
rgb[9401] = 24'b010011101010001111100011;
rgb[9402] = 24'b011010111011001011101000;
rgb[9403] = 24'b100010011100001011101100;
rgb[9404] = 24'b101001101101000111110001;
rgb[9405] = 24'b110001001110000011110101;
rgb[9406] = 24'b111000011110111111111010;
rgb[9407] = 24'b111111111111111111111111;
rgb[9408] = 24'b000000000000000000000000;
rgb[9409] = 24'b000000110001001000011110;
rgb[9410] = 24'b000001100010010100111101;
rgb[9411] = 24'b000010100011100001011011;
rgb[9412] = 24'b000011010100101101111010;
rgb[9413] = 24'b000100000101111010011001;
rgb[9414] = 24'b000101000111000110110111;
rgb[9415] = 24'b000101111000010011010110;
rgb[9416] = 24'b001010001001010111100111;
rgb[9417] = 24'b010001111010010011101010;
rgb[9418] = 24'b011001011011001111101110;
rgb[9419] = 24'b100001001100001011110001;
rgb[9420] = 24'b101000111101000111110100;
rgb[9421] = 24'b110000011110000011111000;
rgb[9422] = 24'b111000001110111111111011;
rgb[9423] = 24'b111111111111111111111111;
rgb[9424] = 24'b000000000000000000000000;
rgb[9425] = 24'b000000100001001100011111;
rgb[9426] = 24'b000001000010011000111111;
rgb[9427] = 24'b000001100011100101011111;
rgb[9428] = 24'b000010010100110001111110;
rgb[9429] = 24'b000010110101111110011110;
rgb[9430] = 24'b000011010111001010111110;
rgb[9431] = 24'b000011111000010111011110;
rgb[9432] = 24'b001000001001011011101111;
rgb[9433] = 24'b010000001010010111110001;
rgb[9434] = 24'b011000001011010011110011;
rgb[9435] = 24'b100000001100001111110101;
rgb[9436] = 24'b100111111101001011111000;
rgb[9437] = 24'b101111111110000111111010;
rgb[9438] = 24'b110111111111000011111100;
rgb[9439] = 24'b111111111111111111111111;
rgb[9440] = 24'b000000000000000000000000;
rgb[9441] = 24'b000000010001001100100000;
rgb[9442] = 24'b000000100010011001000001;
rgb[9443] = 24'b000000110011100101100010;
rgb[9444] = 24'b000001000100110110000011;
rgb[9445] = 24'b000001010110000010100100;
rgb[9446] = 24'b000001100111001111000101;
rgb[9447] = 24'b000001111000011011100110;
rgb[9448] = 24'b000110001001011111110111;
rgb[9449] = 24'b001110011010011011111000;
rgb[9450] = 24'b010110101011010111111001;
rgb[9451] = 24'b011110111100010011111010;
rgb[9452] = 24'b100111001101001011111011;
rgb[9453] = 24'b101111011110000111111100;
rgb[9454] = 24'b110111101111000011111101;
rgb[9455] = 24'b111111111111111111111111;
rgb[9456] = 24'b000000000000000000000000;
rgb[9457] = 24'b000000000001001100100010;
rgb[9458] = 24'b000000000010011001000100;
rgb[9459] = 24'b000000000011101001100110;
rgb[9460] = 24'b000000000100110110001000;
rgb[9461] = 24'b000000000110000110101010;
rgb[9462] = 24'b000000000111010011001100;
rgb[9463] = 24'b000000001000100011101110;
rgb[9464] = 24'b000100011001100111111110;
rgb[9465] = 24'b001100101010011111111111;
rgb[9466] = 24'b010101011011011011111110;
rgb[9467] = 24'b011101101100010011111111;
rgb[9468] = 24'b100110011101001111111111;
rgb[9469] = 24'b101110111110000111111111;
rgb[9470] = 24'b110111011111000011111111;
rgb[9471] = 24'b111111111111111111111111;
rgb[9472] = 24'b000000000000000000000000;
rgb[9473] = 24'b000100010001000100010001;
rgb[9474] = 24'b001000100010001000100010;
rgb[9475] = 24'b001100110011001100110011;
rgb[9476] = 24'b010001000100010001000100;
rgb[9477] = 24'b010101010101010101010101;
rgb[9478] = 24'b011001100110011001100110;
rgb[9479] = 24'b011101110111011101110111;
rgb[9480] = 24'b100010001000100010001000;
rgb[9481] = 24'b100110011001100110011001;
rgb[9482] = 24'b101010101010101010101010;
rgb[9483] = 24'b101110111011101110111011;
rgb[9484] = 24'b110011001100110011001100;
rgb[9485] = 24'b110111011101110111011101;
rgb[9486] = 24'b111011101110111011101110;
rgb[9487] = 24'b111111111111111111111111;
rgb[9488] = 24'b000000000000000000000000;
rgb[9489] = 24'b000011110001000000010010;
rgb[9490] = 24'b000111110010000100100100;
rgb[9491] = 24'b001011110011001000110110;
rgb[9492] = 24'b001111110100001101001000;
rgb[9493] = 24'b010011110101010001011010;
rgb[9494] = 24'b010111110110010101101100;
rgb[9495] = 24'b011011110111011001111110;
rgb[9496] = 24'b100000001000011110001111;
rgb[9497] = 24'b100100101001100010011111;
rgb[9498] = 24'b101001001010100110101111;
rgb[9499] = 24'b101101101011101010111111;
rgb[9500] = 24'b110010001100101111001111;
rgb[9501] = 24'b110110101101110011011111;
rgb[9502] = 24'b111011001110110111101111;
rgb[9503] = 24'b111111111111111111111111;
rgb[9504] = 24'b000000000000000000000000;
rgb[9505] = 24'b000011100001000000010011;
rgb[9506] = 24'b000111010010000100100110;
rgb[9507] = 24'b001011000011001000111001;
rgb[9508] = 24'b001110100100001101001101;
rgb[9509] = 24'b010010010101010001100000;
rgb[9510] = 24'b010110000110010101110011;
rgb[9511] = 24'b011001110111011010000110;
rgb[9512] = 24'b011110001000011110010111;
rgb[9513] = 24'b100010111001100010100110;
rgb[9514] = 24'b100111101010100110110101;
rgb[9515] = 24'b101100011011101011000100;
rgb[9516] = 24'b110001011100101111010010;
rgb[9517] = 24'b110110001101110011100001;
rgb[9518] = 24'b111010111110110111110000;
rgb[9519] = 24'b111111111111111111111111;
rgb[9520] = 24'b000000000000000000000000;
rgb[9521] = 24'b000011010001000000010100;
rgb[9522] = 24'b000110110010000100101000;
rgb[9523] = 24'b001010000011001000111101;
rgb[9524] = 24'b001101100100001101010001;
rgb[9525] = 24'b010001000101010001100101;
rgb[9526] = 24'b010100010110010101111010;
rgb[9527] = 24'b010111110111010110001110;
rgb[9528] = 24'b011100001000011010011111;
rgb[9529] = 24'b100001001001100010101101;
rgb[9530] = 24'b100110001010100110111011;
rgb[9531] = 24'b101011011011101011001000;
rgb[9532] = 24'b110000011100101111010110;
rgb[9533] = 24'b110101101101110011100011;
rgb[9534] = 24'b111010101110110111110001;
rgb[9535] = 24'b111111111111111111111111;
rgb[9536] = 24'b000000000000000000000000;
rgb[9537] = 24'b000011000001000000010101;
rgb[9538] = 24'b000110000010000100101011;
rgb[9539] = 24'b001001010011001001000000;
rgb[9540] = 24'b001100010100001101010110;
rgb[9541] = 24'b001111100101001101101011;
rgb[9542] = 24'b010010100110010010000001;
rgb[9543] = 24'b010101110111010110010110;
rgb[9544] = 24'b011010001000011010100111;
rgb[9545] = 24'b011111011001011110110100;
rgb[9546] = 24'b100100111010100011000000;
rgb[9547] = 24'b101010001011101011001101;
rgb[9548] = 24'b101111101100101111011001;
rgb[9549] = 24'b110100111101110011100110;
rgb[9550] = 24'b111010011110110111110010;
rgb[9551] = 24'b111111111111111111111111;
rgb[9552] = 24'b000000000000000000000000;
rgb[9553] = 24'b000010110001000000010110;
rgb[9554] = 24'b000101100010000100101101;
rgb[9555] = 24'b001000100011001001000100;
rgb[9556] = 24'b001011010100001001011010;
rgb[9557] = 24'b001110000101001101110001;
rgb[9558] = 24'b010001000110010010001000;
rgb[9559] = 24'b010011110111010110011110;
rgb[9560] = 24'b011000001000011010101111;
rgb[9561] = 24'b011101101001011110111011;
rgb[9562] = 24'b100011011010100011000110;
rgb[9563] = 24'b101001001011100111010001;
rgb[9564] = 24'b101110111100101111011101;
rgb[9565] = 24'b110100011101110011101000;
rgb[9566] = 24'b111010001110110111110011;
rgb[9567] = 24'b111111111111111111111111;
rgb[9568] = 24'b000000000000000000000000;
rgb[9569] = 24'b000010100001000000010111;
rgb[9570] = 24'b000101000010000100101111;
rgb[9571] = 24'b000111100011001001000111;
rgb[9572] = 24'b001010000100001001011111;
rgb[9573] = 24'b001100110101001101110110;
rgb[9574] = 24'b001111010110010010001110;
rgb[9575] = 24'b010001110111010010100110;
rgb[9576] = 24'b010110001000010110110111;
rgb[9577] = 24'b011100001001011111000001;
rgb[9578] = 24'b100001111010100011001100;
rgb[9579] = 24'b100111111011100111010110;
rgb[9580] = 24'b101101111100101111100000;
rgb[9581] = 24'b110011111101110011101010;
rgb[9582] = 24'b111001111110110111110100;
rgb[9583] = 24'b111111111111111111111110;
rgb[9584] = 24'b000000000000000000000000;
rgb[9585] = 24'b000010010001000000011000;
rgb[9586] = 24'b000100100010000100110001;
rgb[9587] = 24'b000110110011000101001010;
rgb[9588] = 24'b001001000100001001100011;
rgb[9589] = 24'b001011010101001101111100;
rgb[9590] = 24'b001101100110001110010101;
rgb[9591] = 24'b001111110111010010101110;
rgb[9592] = 24'b010100001000010110111111;
rgb[9593] = 24'b011010011001011011001000;
rgb[9594] = 24'b100000101010100011010001;
rgb[9595] = 24'b100110111011100111011010;
rgb[9596] = 24'b101101001100101011100011;
rgb[9597] = 24'b110011011101110011101100;
rgb[9598] = 24'b111001101110110111110101;
rgb[9599] = 24'b111111111111111111111111;
rgb[9600] = 24'b000000000000000000000000;
rgb[9601] = 24'b000001110001000000011010;
rgb[9602] = 24'b000011110010000100110100;
rgb[9603] = 24'b000101110011000101001110;
rgb[9604] = 24'b000111110100001001101000;
rgb[9605] = 24'b001001110101001010000010;
rgb[9606] = 24'b001011110110001110011100;
rgb[9607] = 24'b001101110111001110110110;
rgb[9608] = 24'b010010001000010011000111;
rgb[9609] = 24'b011000101001011011001111;
rgb[9610] = 24'b011111001010011111010111;
rgb[9611] = 24'b100101101011100111011111;
rgb[9612] = 24'b101100001100101011100111;
rgb[9613] = 24'b110010101101110011101111;
rgb[9614] = 24'b111001001110110111110111;
rgb[9615] = 24'b111111111111111111111110;
rgb[9616] = 24'b000000000000000000000000;
rgb[9617] = 24'b000001100001000000011011;
rgb[9618] = 24'b000011010010000100110110;
rgb[9619] = 24'b000101000011000101010001;
rgb[9620] = 24'b000110110100001001101100;
rgb[9621] = 24'b001000010101001010001000;
rgb[9622] = 24'b001010000110001110100011;
rgb[9623] = 24'b001011110111001110111110;
rgb[9624] = 24'b010000001000010011001111;
rgb[9625] = 24'b010110111001011011010110;
rgb[9626] = 24'b011101101010011111011101;
rgb[9627] = 24'b100100101011100111100011;
rgb[9628] = 24'b101011011100101011101010;
rgb[9629] = 24'b110010001101110011110001;
rgb[9630] = 24'b111000111110110111111000;
rgb[9631] = 24'b111111111111111111111111;
rgb[9632] = 24'b000000000000000000000000;
rgb[9633] = 24'b000001010001000000011100;
rgb[9634] = 24'b000010110010000000111000;
rgb[9635] = 24'b000100010011000101010101;
rgb[9636] = 24'b000101100100000101110001;
rgb[9637] = 24'b000111000101001010001101;
rgb[9638] = 24'b001000100110001010101010;
rgb[9639] = 24'b001001110111001111000110;
rgb[9640] = 24'b001110001000010011010111;
rgb[9641] = 24'b010101001001010111011101;
rgb[9642] = 24'b011100011010011111100010;
rgb[9643] = 24'b100011011011100011101000;
rgb[9644] = 24'b101010101100101011101110;
rgb[9645] = 24'b110001101101101111110011;
rgb[9646] = 24'b111000101110110111111001;
rgb[9647] = 24'b111111111111111111111110;
rgb[9648] = 24'b000000000000000000000000;
rgb[9649] = 24'b000001000001000000011101;
rgb[9650] = 24'b000010010010000000111010;
rgb[9651] = 24'b000011010011000101011000;
rgb[9652] = 24'b000100100100000101110101;
rgb[9653] = 24'b000101100101001010010011;
rgb[9654] = 24'b000110110110001010110000;
rgb[9655] = 24'b000111110111001011001110;
rgb[9656] = 24'b001100001000001111011111;
rgb[9657] = 24'b010011101001010111100011;
rgb[9658] = 24'b011010111010011111101000;
rgb[9659] = 24'b100010011011100011101100;
rgb[9660] = 24'b101001101100101011110001;
rgb[9661] = 24'b110001001101101111110101;
rgb[9662] = 24'b111000011110110111111010;
rgb[9663] = 24'b111111111111111111111111;
rgb[9664] = 24'b000000000000000000000000;
rgb[9665] = 24'b000000110001000000011110;
rgb[9666] = 24'b000001100010000000111101;
rgb[9667] = 24'b000010100011000101011011;
rgb[9668] = 24'b000011010100000101111010;
rgb[9669] = 24'b000100000101000110011001;
rgb[9670] = 24'b000101000110001010110111;
rgb[9671] = 24'b000101110111001011010110;
rgb[9672] = 24'b001010001000001111100111;
rgb[9673] = 24'b010001111001010111101010;
rgb[9674] = 24'b011001011010011011101110;
rgb[9675] = 24'b100001001011100011110001;
rgb[9676] = 24'b101000111100101011110100;
rgb[9677] = 24'b110000011101101111111000;
rgb[9678] = 24'b111000001110110111111011;
rgb[9679] = 24'b111111111111111111111111;
rgb[9680] = 24'b000000000000000000000000;
rgb[9681] = 24'b000000100001000000011111;
rgb[9682] = 24'b000001000010000000111111;
rgb[9683] = 24'b000001100011000001011111;
rgb[9684] = 24'b000010010100000101111110;
rgb[9685] = 24'b000010110101000110011110;
rgb[9686] = 24'b000011010110000110111110;
rgb[9687] = 24'b000011110111001011011110;
rgb[9688] = 24'b001000001000001111101111;
rgb[9689] = 24'b010000001001010011110001;
rgb[9690] = 24'b011000001010011011110011;
rgb[9691] = 24'b100000001011100011110101;
rgb[9692] = 24'b100111111100100111111000;
rgb[9693] = 24'b101111111101101111111010;
rgb[9694] = 24'b110111111110110111111100;
rgb[9695] = 24'b111111111111111111111111;
rgb[9696] = 24'b000000000000000000000000;
rgb[9697] = 24'b000000010001000000100000;
rgb[9698] = 24'b000000100010000001000001;
rgb[9699] = 24'b000000110011000001100010;
rgb[9700] = 24'b000001000100000010000011;
rgb[9701] = 24'b000001010101000110100100;
rgb[9702] = 24'b000001100110000111000101;
rgb[9703] = 24'b000001110111000111100110;
rgb[9704] = 24'b000110001000001011110111;
rgb[9705] = 24'b001110011001010011111000;
rgb[9706] = 24'b010110101010011011111001;
rgb[9707] = 24'b011110111011011111111010;
rgb[9708] = 24'b100111001100100111111011;
rgb[9709] = 24'b101111011101101111111100;
rgb[9710] = 24'b110111101110110111111101;
rgb[9711] = 24'b111111111111111111111111;
rgb[9712] = 24'b000000000000000000000000;
rgb[9713] = 24'b000000000001000000100010;
rgb[9714] = 24'b000000000010000001000100;
rgb[9715] = 24'b000000000011000001100110;
rgb[9716] = 24'b000000000100000010001000;
rgb[9717] = 24'b000000000101000010101010;
rgb[9718] = 24'b000000000110000111001100;
rgb[9719] = 24'b000000000111000111101110;
rgb[9720] = 24'b000100011000001011111110;
rgb[9721] = 24'b001100101001010011111111;
rgb[9722] = 24'b010101011010010111111110;
rgb[9723] = 24'b011101101011011111111111;
rgb[9724] = 24'b100110011100100111111111;
rgb[9725] = 24'b101110111101101111111111;
rgb[9726] = 24'b110111011110110111111111;
rgb[9727] = 24'b111111111111111111111111;
rgb[9728] = 24'b000000000000000000000000;
rgb[9729] = 24'b000100010001000100010001;
rgb[9730] = 24'b001000100010001000100010;
rgb[9731] = 24'b001100110011001100110011;
rgb[9732] = 24'b010001000100010001000100;
rgb[9733] = 24'b010101010101010101010101;
rgb[9734] = 24'b011001100110011001100110;
rgb[9735] = 24'b011101110111011101110111;
rgb[9736] = 24'b100010001000100010001000;
rgb[9737] = 24'b100110011001100110011001;
rgb[9738] = 24'b101010101010101010101010;
rgb[9739] = 24'b101110111011101110111011;
rgb[9740] = 24'b110011001100110011001100;
rgb[9741] = 24'b110111011101110111011101;
rgb[9742] = 24'b111011101110111011101110;
rgb[9743] = 24'b111111111111111111111111;
rgb[9744] = 24'b000000000000000000000000;
rgb[9745] = 24'b000011110001000000010010;
rgb[9746] = 24'b000111110010000100100100;
rgb[9747] = 24'b001011110011001000110110;
rgb[9748] = 24'b001111110100001001001000;
rgb[9749] = 24'b010011110101001101011010;
rgb[9750] = 24'b010111110110010001101100;
rgb[9751] = 24'b011011110111010101111110;
rgb[9752] = 24'b100000001000011010001111;
rgb[9753] = 24'b100100101001011110011111;
rgb[9754] = 24'b101001001010100010101111;
rgb[9755] = 24'b101101101011100110111111;
rgb[9756] = 24'b110010001100101111001111;
rgb[9757] = 24'b110110101101110011011111;
rgb[9758] = 24'b111011001110110111101111;
rgb[9759] = 24'b111111111111111111111111;
rgb[9760] = 24'b000000000000000000000000;
rgb[9761] = 24'b000011100001000000010011;
rgb[9762] = 24'b000111010010000000100110;
rgb[9763] = 24'b001011000011000100111001;
rgb[9764] = 24'b001110100100000101001101;
rgb[9765] = 24'b010010010101001001100000;
rgb[9766] = 24'b010110000110001001110011;
rgb[9767] = 24'b011001110111001110000110;
rgb[9768] = 24'b011110001000010010010111;
rgb[9769] = 24'b100010111001010110100110;
rgb[9770] = 24'b100111101010011110110101;
rgb[9771] = 24'b101100011011100011000100;
rgb[9772] = 24'b110001011100101011010010;
rgb[9773] = 24'b110110001101101111100001;
rgb[9774] = 24'b111010111110110111110000;
rgb[9775] = 24'b111111111111111111111111;
rgb[9776] = 24'b000000000000000000000000;
rgb[9777] = 24'b000011010001000000010100;
rgb[9778] = 24'b000110110010000000101000;
rgb[9779] = 24'b001010000011000000111101;
rgb[9780] = 24'b001101100100000001010001;
rgb[9781] = 24'b010001000101000001100101;
rgb[9782] = 24'b010100010110000101111010;
rgb[9783] = 24'b010111110111000110001110;
rgb[9784] = 24'b011100001000001010011111;
rgb[9785] = 24'b100001001001010010101101;
rgb[9786] = 24'b100110001010010110111011;
rgb[9787] = 24'b101011011011011111001000;
rgb[9788] = 24'b110000011100100111010110;
rgb[9789] = 24'b110101101101101111100011;
rgb[9790] = 24'b111010101110110111110001;
rgb[9791] = 24'b111111111111111111111111;
rgb[9792] = 24'b000000000000000000000000;
rgb[9793] = 24'b000011000000111100010101;
rgb[9794] = 24'b000110000001111100101011;
rgb[9795] = 24'b001001010010111101000000;
rgb[9796] = 24'b001100010011111101010110;
rgb[9797] = 24'b001111100100111101101011;
rgb[9798] = 24'b010010100101111110000001;
rgb[9799] = 24'b010101110110111110010110;
rgb[9800] = 24'b011010001000000010100111;
rgb[9801] = 24'b011111011001001010110100;
rgb[9802] = 24'b100100111010010011000000;
rgb[9803] = 24'b101010001011011011001101;
rgb[9804] = 24'b101111101100100011011001;
rgb[9805] = 24'b110100111101101011100110;
rgb[9806] = 24'b111010011110110011110010;
rgb[9807] = 24'b111111111111111111111111;
rgb[9808] = 24'b000000000000000000000000;
rgb[9809] = 24'b000010110000111100010110;
rgb[9810] = 24'b000101100001111100101101;
rgb[9811] = 24'b001000100010111001000100;
rgb[9812] = 24'b001011010011111001011010;
rgb[9813] = 24'b001110000100111001110001;
rgb[9814] = 24'b010001000101110110001000;
rgb[9815] = 24'b010011110110110110011110;
rgb[9816] = 24'b011000000111111010101111;
rgb[9817] = 24'b011101101001000010111011;
rgb[9818] = 24'b100011011010001111000110;
rgb[9819] = 24'b101001001011010111010001;
rgb[9820] = 24'b101110111100011111011101;
rgb[9821] = 24'b110100011101101011101000;
rgb[9822] = 24'b111010001110110011110011;
rgb[9823] = 24'b111111111111111111111111;
rgb[9824] = 24'b000000000000000000000000;
rgb[9825] = 24'b000010100000111100010111;
rgb[9826] = 24'b000101000001111000101111;
rgb[9827] = 24'b000111100010111001000111;
rgb[9828] = 24'b001010000011110101011111;
rgb[9829] = 24'b001100110100110001110110;
rgb[9830] = 24'b001111010101110010001110;
rgb[9831] = 24'b010001110110101110100110;
rgb[9832] = 24'b010110000111110010110111;
rgb[9833] = 24'b011100001000111111000001;
rgb[9834] = 24'b100001111010000111001100;
rgb[9835] = 24'b100111111011010011010110;
rgb[9836] = 24'b101101111100011111100000;
rgb[9837] = 24'b110011111101100111101010;
rgb[9838] = 24'b111001111110110011110100;
rgb[9839] = 24'b111111111111111111111110;
rgb[9840] = 24'b000000000000000000000000;
rgb[9841] = 24'b000010010000111100011000;
rgb[9842] = 24'b000100100001111000110001;
rgb[9843] = 24'b000110110010110101001010;
rgb[9844] = 24'b001001000011110001100011;
rgb[9845] = 24'b001011010100101101111100;
rgb[9846] = 24'b001101100101101010010101;
rgb[9847] = 24'b001111110110100110101110;
rgb[9848] = 24'b010100000111101010111111;
rgb[9849] = 24'b011010011000110111001000;
rgb[9850] = 24'b100000101010000011010001;
rgb[9851] = 24'b100110111011001111011010;
rgb[9852] = 24'b101101001100011011100011;
rgb[9853] = 24'b110011011101100111101100;
rgb[9854] = 24'b111001101110110011110101;
rgb[9855] = 24'b111111111111111111111111;
rgb[9856] = 24'b000000000000000000000000;
rgb[9857] = 24'b000001110000111000011010;
rgb[9858] = 24'b000011110001110100110100;
rgb[9859] = 24'b000101110010110001001110;
rgb[9860] = 24'b000111110011101101101000;
rgb[9861] = 24'b001001110100101010000010;
rgb[9862] = 24'b001011110101100110011100;
rgb[9863] = 24'b001101110110011110110110;
rgb[9864] = 24'b010010000111100011000111;
rgb[9865] = 24'b011000101000110011001111;
rgb[9866] = 24'b011111001001111111010111;
rgb[9867] = 24'b100101101011001011011111;
rgb[9868] = 24'b101100001100010111100111;
rgb[9869] = 24'b110010101101100011101111;
rgb[9870] = 24'b111001001110101111110111;
rgb[9871] = 24'b111111111111111111111110;
rgb[9872] = 24'b000000000000000000000000;
rgb[9873] = 24'b000001100000111000011011;
rgb[9874] = 24'b000011010001110100110110;
rgb[9875] = 24'b000101000010101101010001;
rgb[9876] = 24'b000110110011101001101100;
rgb[9877] = 24'b001000010100100010001000;
rgb[9878] = 24'b001010000101011110100011;
rgb[9879] = 24'b001011110110010110111110;
rgb[9880] = 24'b010000000111011111001111;
rgb[9881] = 24'b010110111000101011010110;
rgb[9882] = 24'b011101101001110111011101;
rgb[9883] = 24'b100100101011000111100011;
rgb[9884] = 24'b101011011100010011101010;
rgb[9885] = 24'b110010001101100011110001;
rgb[9886] = 24'b111000111110101111111000;
rgb[9887] = 24'b111111111111111111111111;
rgb[9888] = 24'b000000000000000000000000;
rgb[9889] = 24'b000001010000111000011100;
rgb[9890] = 24'b000010110001110000111000;
rgb[9891] = 24'b000100010010101001010101;
rgb[9892] = 24'b000101100011100101110001;
rgb[9893] = 24'b000111000100011110001101;
rgb[9894] = 24'b001000100101010110101010;
rgb[9895] = 24'b001001110110010011000110;
rgb[9896] = 24'b001110000111010111010111;
rgb[9897] = 24'b010101001000100011011101;
rgb[9898] = 24'b011100011001110011100010;
rgb[9899] = 24'b100011011011000011101000;
rgb[9900] = 24'b101010101100001111101110;
rgb[9901] = 24'b110001101101011111110011;
rgb[9902] = 24'b111000101110101111111001;
rgb[9903] = 24'b111111111111111111111110;
rgb[9904] = 24'b000000000000000000000000;
rgb[9905] = 24'b000001000000111000011101;
rgb[9906] = 24'b000010010001110000111010;
rgb[9907] = 24'b000011010010101001011000;
rgb[9908] = 24'b000100100011100001110101;
rgb[9909] = 24'b000101100100011010010011;
rgb[9910] = 24'b000110110101010010110000;
rgb[9911] = 24'b000111110110001011001110;
rgb[9912] = 24'b001100000111001111011111;
rgb[9913] = 24'b010011101000011111100011;
rgb[9914] = 24'b011010111001101111101000;
rgb[9915] = 24'b100010011010111111101100;
rgb[9916] = 24'b101001101100001111110001;
rgb[9917] = 24'b110001001101011111110101;
rgb[9918] = 24'b111000011110101111111010;
rgb[9919] = 24'b111111111111111111111111;
rgb[9920] = 24'b000000000000000000000000;
rgb[9921] = 24'b000000110000110100011110;
rgb[9922] = 24'b000001100001101100111101;
rgb[9923] = 24'b000010100010100101011011;
rgb[9924] = 24'b000011010011011101111010;
rgb[9925] = 24'b000100000100010010011001;
rgb[9926] = 24'b000101000101001010110111;
rgb[9927] = 24'b000101110110000011010110;
rgb[9928] = 24'b001010000111000111100111;
rgb[9929] = 24'b010001111000010111101010;
rgb[9930] = 24'b011001011001100111101110;
rgb[9931] = 24'b100001001010111011110001;
rgb[9932] = 24'b101000111100001011110100;
rgb[9933] = 24'b110000011101011011111000;
rgb[9934] = 24'b111000001110101011111011;
rgb[9935] = 24'b111111111111111111111111;
rgb[9936] = 24'b000000000000000000000000;
rgb[9937] = 24'b000000100000110100011111;
rgb[9938] = 24'b000001000001101000111111;
rgb[9939] = 24'b000001100010100001011111;
rgb[9940] = 24'b000010010011010101111110;
rgb[9941] = 24'b000010110100001110011110;
rgb[9942] = 24'b000011010101000010111110;
rgb[9943] = 24'b000011110101111011011110;
rgb[9944] = 24'b001000000110111111101111;
rgb[9945] = 24'b010000001000001111110001;
rgb[9946] = 24'b011000001001100011110011;
rgb[9947] = 24'b100000001010110011110101;
rgb[9948] = 24'b100111111100000111111000;
rgb[9949] = 24'b101111111101010111111010;
rgb[9950] = 24'b110111111110101011111100;
rgb[9951] = 24'b111111111111111111111111;
rgb[9952] = 24'b000000000000000000000000;
rgb[9953] = 24'b000000010000110100100000;
rgb[9954] = 24'b000000100001101001000001;
rgb[9955] = 24'b000000110010011101100010;
rgb[9956] = 24'b000001000011010010000011;
rgb[9957] = 24'b000001010100001010100100;
rgb[9958] = 24'b000001100100111111000101;
rgb[9959] = 24'b000001110101110011100110;
rgb[9960] = 24'b000110000110110111110111;
rgb[9961] = 24'b001110011000001011111000;
rgb[9962] = 24'b010110101001011111111001;
rgb[9963] = 24'b011110111010101111111010;
rgb[9964] = 24'b100111001100000011111011;
rgb[9965] = 24'b101111011101010111111100;
rgb[9966] = 24'b110111101110101011111101;
rgb[9967] = 24'b111111111111111111111111;
rgb[9968] = 24'b000000000000000000000000;
rgb[9969] = 24'b000000000000110000100010;
rgb[9970] = 24'b000000000001100101000100;
rgb[9971] = 24'b000000000010011001100110;
rgb[9972] = 24'b000000000011001110001000;
rgb[9973] = 24'b000000000100000010101010;
rgb[9974] = 24'b000000000100110111001100;
rgb[9975] = 24'b000000000101101011101110;
rgb[9976] = 24'b000100010110101111111110;
rgb[9977] = 24'b001100101000000011111111;
rgb[9978] = 24'b010101011001010111111110;
rgb[9979] = 24'b011101101010101011111111;
rgb[9980] = 24'b100110011011111111111111;
rgb[9981] = 24'b101110111101010011111111;
rgb[9982] = 24'b110111011110100111111111;
rgb[9983] = 24'b111111111111111111111111;
rgb[9984] = 24'b000000000000000000000000;
rgb[9985] = 24'b000100010001000100010001;
rgb[9986] = 24'b001000100010001000100010;
rgb[9987] = 24'b001100110011001100110011;
rgb[9988] = 24'b010001000100010001000100;
rgb[9989] = 24'b010101010101010101010101;
rgb[9990] = 24'b011001100110011001100110;
rgb[9991] = 24'b011101110111011101110111;
rgb[9992] = 24'b100010001000100010001000;
rgb[9993] = 24'b100110011001100110011001;
rgb[9994] = 24'b101010101010101010101010;
rgb[9995] = 24'b101110111011101110111011;
rgb[9996] = 24'b110011001100110011001100;
rgb[9997] = 24'b110111011101110111011101;
rgb[9998] = 24'b111011101110111011101110;
rgb[9999] = 24'b111111111111111111111111;
rgb[10000] = 24'b000000000000000000000000;
rgb[10001] = 24'b000011110001000000010010;
rgb[10002] = 24'b000111110010000100100100;
rgb[10003] = 24'b001011110011000100110110;
rgb[10004] = 24'b001111110100001001001000;
rgb[10005] = 24'b010011110101001001011010;
rgb[10006] = 24'b010111110110001101101100;
rgb[10007] = 24'b011011110111001101111110;
rgb[10008] = 24'b100000001000010010001111;
rgb[10009] = 24'b100100101001011010011111;
rgb[10010] = 24'b101001001010011110101111;
rgb[10011] = 24'b101101101011100110111111;
rgb[10012] = 24'b110010001100101011001111;
rgb[10013] = 24'b110110101101110011011111;
rgb[10014] = 24'b111011001110110111101111;
rgb[10015] = 24'b111111111111111111111111;
rgb[10016] = 24'b000000000000000000000000;
rgb[10017] = 24'b000011100001000000010011;
rgb[10018] = 24'b000111010010000000100110;
rgb[10019] = 24'b001011000011000000111001;
rgb[10020] = 24'b001110100100000001001101;
rgb[10021] = 24'b010010010101000001100000;
rgb[10022] = 24'b010110000110000001110011;
rgb[10023] = 24'b011001110111000010000110;
rgb[10024] = 24'b011110001000000110010111;
rgb[10025] = 24'b100010111001001110100110;
rgb[10026] = 24'b100111101010010110110101;
rgb[10027] = 24'b101100011011011111000100;
rgb[10028] = 24'b110001011100100111010010;
rgb[10029] = 24'b110110001101101111100001;
rgb[10030] = 24'b111010111110110111110000;
rgb[10031] = 24'b111111111111111111111111;
rgb[10032] = 24'b000000000000000000000000;
rgb[10033] = 24'b000011010000111100010100;
rgb[10034] = 24'b000110110001111100101000;
rgb[10035] = 24'b001010000010111000111101;
rgb[10036] = 24'b001101100011111001010001;
rgb[10037] = 24'b010001000100110101100101;
rgb[10038] = 24'b010100010101110101111010;
rgb[10039] = 24'b010111110110110010001110;
rgb[10040] = 24'b011100000111110110011111;
rgb[10041] = 24'b100001001001000010101101;
rgb[10042] = 24'b100110001010001010111011;
rgb[10043] = 24'b101011011011010111001000;
rgb[10044] = 24'b110000011100011111010110;
rgb[10045] = 24'b110101101101101011100011;
rgb[10046] = 24'b111010101110110011110001;
rgb[10047] = 24'b111111111111111111111111;
rgb[10048] = 24'b000000000000000000000000;
rgb[10049] = 24'b000011000000111100010101;
rgb[10050] = 24'b000110000001111000101011;
rgb[10051] = 24'b001001010010110101000000;
rgb[10052] = 24'b001100010011110001010110;
rgb[10053] = 24'b001111100100101101101011;
rgb[10054] = 24'b010010100101101010000001;
rgb[10055] = 24'b010101110110100110010110;
rgb[10056] = 24'b011010000111101010100111;
rgb[10057] = 24'b011111011000110110110100;
rgb[10058] = 24'b100100111010000011000000;
rgb[10059] = 24'b101010001011001111001101;
rgb[10060] = 24'b101111101100011011011001;
rgb[10061] = 24'b110100111101100111100110;
rgb[10062] = 24'b111010011110110011110010;
rgb[10063] = 24'b111111111111111111111111;
rgb[10064] = 24'b000000000000000000000000;
rgb[10065] = 24'b000010110000111000010110;
rgb[10066] = 24'b000101100001110100101101;
rgb[10067] = 24'b001000100010101101000100;
rgb[10068] = 24'b001011010011101001011010;
rgb[10069] = 24'b001110000100100001110001;
rgb[10070] = 24'b010001000101011110001000;
rgb[10071] = 24'b010011110110010110011110;
rgb[10072] = 24'b011000000111011010101111;
rgb[10073] = 24'b011101101000101010111011;
rgb[10074] = 24'b100011011001110111000110;
rgb[10075] = 24'b101001001011000111010001;
rgb[10076] = 24'b101110111100010011011101;
rgb[10077] = 24'b110100011101100011101000;
rgb[10078] = 24'b111010001110101111110011;
rgb[10079] = 24'b111111111111111111111111;
rgb[10080] = 24'b000000000000000000000000;
rgb[10081] = 24'b000010100000111000010111;
rgb[10082] = 24'b000101000001110000101111;
rgb[10083] = 24'b000111100010101001000111;
rgb[10084] = 24'b001010000011100001011111;
rgb[10085] = 24'b001100110100011001110110;
rgb[10086] = 24'b001111010101010010001110;
rgb[10087] = 24'b010001110110001010100110;
rgb[10088] = 24'b010110000111001110110111;
rgb[10089] = 24'b011100001000011111000001;
rgb[10090] = 24'b100001111001101111001100;
rgb[10091] = 24'b100111111010111111010110;
rgb[10092] = 24'b101101111100001111100000;
rgb[10093] = 24'b110011111101011111101010;
rgb[10094] = 24'b111001111110101111110100;
rgb[10095] = 24'b111111111111111111111110;
rgb[10096] = 24'b000000000000000000000000;
rgb[10097] = 24'b000010010000110100011000;
rgb[10098] = 24'b000100100001101100110001;
rgb[10099] = 24'b000110110010100001001010;
rgb[10100] = 24'b001001000011011001100011;
rgb[10101] = 24'b001011010100001101111100;
rgb[10102] = 24'b001101100101000110010101;
rgb[10103] = 24'b001111110101111110101110;
rgb[10104] = 24'b010100000111000010111111;
rgb[10105] = 24'b011010011000010011001000;
rgb[10106] = 24'b100000101001100011010001;
rgb[10107] = 24'b100110111010110111011010;
rgb[10108] = 24'b101101001100000111100011;
rgb[10109] = 24'b110011011101011011101100;
rgb[10110] = 24'b111001101110101011110101;
rgb[10111] = 24'b111111111111111111111111;
rgb[10112] = 24'b000000000000000000000000;
rgb[10113] = 24'b000001110000110100011010;
rgb[10114] = 24'b000011110001101000110100;
rgb[10115] = 24'b000101110010011101001110;
rgb[10116] = 24'b000111110011010001101000;
rgb[10117] = 24'b001001110100000110000010;
rgb[10118] = 24'b001011110100111010011100;
rgb[10119] = 24'b001101110101101110110110;
rgb[10120] = 24'b010010000110110011000111;
rgb[10121] = 24'b011000101000000111001111;
rgb[10122] = 24'b011111001001011011010111;
rgb[10123] = 24'b100101101010101111011111;
rgb[10124] = 24'b101100001100000011100111;
rgb[10125] = 24'b110010101101010111101111;
rgb[10126] = 24'b111001001110101011110111;
rgb[10127] = 24'b111111111111111111111110;
rgb[10128] = 24'b000000000000000000000000;
rgb[10129] = 24'b000001100000110000011011;
rgb[10130] = 24'b000011010001100100110110;
rgb[10131] = 24'b000101000010010101010001;
rgb[10132] = 24'b000110110011001001101100;
rgb[10133] = 24'b001000010011111110001000;
rgb[10134] = 24'b001010000100101110100011;
rgb[10135] = 24'b001011110101100010111110;
rgb[10136] = 24'b010000000110100111001111;
rgb[10137] = 24'b010110110111111011010110;
rgb[10138] = 24'b011101101001010011011101;
rgb[10139] = 24'b100100101010100111100011;
rgb[10140] = 24'b101011011011111011101010;
rgb[10141] = 24'b110010001101010011110001;
rgb[10142] = 24'b111000111110100111111000;
rgb[10143] = 24'b111111111111111111111111;
rgb[10144] = 24'b000000000000000000000000;
rgb[10145] = 24'b000001010000110000011100;
rgb[10146] = 24'b000010110001100000111000;
rgb[10147] = 24'b000100010010010001010101;
rgb[10148] = 24'b000101100011000001110001;
rgb[10149] = 24'b000111000011110010001101;
rgb[10150] = 24'b001000100100100010101010;
rgb[10151] = 24'b001001110101010011000110;
rgb[10152] = 24'b001110000110010111010111;
rgb[10153] = 24'b010101000111101111011101;
rgb[10154] = 24'b011100011001000111100010;
rgb[10155] = 24'b100011011010011111101000;
rgb[10156] = 24'b101010101011110111101110;
rgb[10157] = 24'b110001101101001111110011;
rgb[10158] = 24'b111000101110100111111001;
rgb[10159] = 24'b111111111111111111111110;
rgb[10160] = 24'b000000000000000000000000;
rgb[10161] = 24'b000001000000101100011101;
rgb[10162] = 24'b000010010001011100111010;
rgb[10163] = 24'b000011010010001001011000;
rgb[10164] = 24'b000100100010111001110101;
rgb[10165] = 24'b000101100011101010010011;
rgb[10166] = 24'b000110110100010110110000;
rgb[10167] = 24'b000111110101000111001110;
rgb[10168] = 24'b001100000110001011011111;
rgb[10169] = 24'b010011100111100011100011;
rgb[10170] = 24'b011010111000111111101000;
rgb[10171] = 24'b100010011010010111101100;
rgb[10172] = 24'b101001101011101111110001;
rgb[10173] = 24'b110001001101001011110101;
rgb[10174] = 24'b111000011110100011111010;
rgb[10175] = 24'b111111111111111111111111;
rgb[10176] = 24'b000000000000000000000000;
rgb[10177] = 24'b000000110000101100011110;
rgb[10178] = 24'b000001100001011000111101;
rgb[10179] = 24'b000010100010000101011011;
rgb[10180] = 24'b000011010010110001111010;
rgb[10181] = 24'b000100000011011110011001;
rgb[10182] = 24'b000101000100001110110111;
rgb[10183] = 24'b000101110100111011010110;
rgb[10184] = 24'b001010000101111111100111;
rgb[10185] = 24'b010001110111011011101010;
rgb[10186] = 24'b011001011000110011101110;
rgb[10187] = 24'b100001001010001111110001;
rgb[10188] = 24'b101000111011101011110100;
rgb[10189] = 24'b110000011101000111111000;
rgb[10190] = 24'b111000001110100011111011;
rgb[10191] = 24'b111111111111111111111111;
rgb[10192] = 24'b000000000000000000000000;
rgb[10193] = 24'b000000100000101000011111;
rgb[10194] = 24'b000001000001010100111111;
rgb[10195] = 24'b000001100010000001011111;
rgb[10196] = 24'b000010010010101001111110;
rgb[10197] = 24'b000010110011010110011110;
rgb[10198] = 24'b000011010100000010111110;
rgb[10199] = 24'b000011110100101011011110;
rgb[10200] = 24'b001000000101101111101111;
rgb[10201] = 24'b010000000111001111110001;
rgb[10202] = 24'b011000001000101011110011;
rgb[10203] = 24'b100000001010000111110101;
rgb[10204] = 24'b100111111011100111111000;
rgb[10205] = 24'b101111111101000011111010;
rgb[10206] = 24'b110111111110011111111100;
rgb[10207] = 24'b111111111111111111111111;
rgb[10208] = 24'b000000000000000000000000;
rgb[10209] = 24'b000000010000101000100000;
rgb[10210] = 24'b000000100001010001000001;
rgb[10211] = 24'b000000110001111001100010;
rgb[10212] = 24'b000001000010100010000011;
rgb[10213] = 24'b000001010011001010100100;
rgb[10214] = 24'b000001100011110111000101;
rgb[10215] = 24'b000001110100011111100110;
rgb[10216] = 24'b000110000101100011110111;
rgb[10217] = 24'b001110010111000011111000;
rgb[10218] = 24'b010110101000011111111001;
rgb[10219] = 24'b011110111001111111111010;
rgb[10220] = 24'b100111001011011111111011;
rgb[10221] = 24'b101111011100111111111100;
rgb[10222] = 24'b110111101110011111111101;
rgb[10223] = 24'b111111111111111111111111;
rgb[10224] = 24'b000000000000000000000000;
rgb[10225] = 24'b000000000000100100100010;
rgb[10226] = 24'b000000000001001101000100;
rgb[10227] = 24'b000000000001110101100110;
rgb[10228] = 24'b000000000010011010001000;
rgb[10229] = 24'b000000000011000010101010;
rgb[10230] = 24'b000000000011101011001100;
rgb[10231] = 24'b000000000100001111101110;
rgb[10232] = 24'b000100010101010011111110;
rgb[10233] = 24'b001100100110110111111111;
rgb[10234] = 24'b010101011000010111111110;
rgb[10235] = 24'b011101101001110111111111;
rgb[10236] = 24'b100110011011011011111111;
rgb[10237] = 24'b101110111100111011111111;
rgb[10238] = 24'b110111011110011011111111;
rgb[10239] = 24'b111111111111111111111111;
rgb[10240] = 24'b000000000000000000000000;
rgb[10241] = 24'b000100010001000100010001;
rgb[10242] = 24'b001000100010001000100010;
rgb[10243] = 24'b001100110011001100110011;
rgb[10244] = 24'b010001000100010001000100;
rgb[10245] = 24'b010101010101010101010101;
rgb[10246] = 24'b011001100110011001100110;
rgb[10247] = 24'b011101110111011101110111;
rgb[10248] = 24'b100010001000100010001000;
rgb[10249] = 24'b100110011001100110011001;
rgb[10250] = 24'b101010101010101010101010;
rgb[10251] = 24'b101110111011101110111011;
rgb[10252] = 24'b110011001100110011001100;
rgb[10253] = 24'b110111011101110111011101;
rgb[10254] = 24'b111011101110111011101110;
rgb[10255] = 24'b111111111111111111111111;
rgb[10256] = 24'b000000000000000000000000;
rgb[10257] = 24'b000011110001000000010010;
rgb[10258] = 24'b000111110010000000100100;
rgb[10259] = 24'b001011110011000000110110;
rgb[10260] = 24'b001111110100000101001000;
rgb[10261] = 24'b010011110101000101011010;
rgb[10262] = 24'b010111110110000101101100;
rgb[10263] = 24'b011011110111001001111110;
rgb[10264] = 24'b100000001000001110001111;
rgb[10265] = 24'b100100101001010010011111;
rgb[10266] = 24'b101001001010011010101111;
rgb[10267] = 24'b101101101011100010111111;
rgb[10268] = 24'b110010001100100111001111;
rgb[10269] = 24'b110110101101101111011111;
rgb[10270] = 24'b111011001110110111101111;
rgb[10271] = 24'b111111111111111111111111;
rgb[10272] = 24'b000000000000000000000000;
rgb[10273] = 24'b000011100000111100010011;
rgb[10274] = 24'b000111010001111100100110;
rgb[10275] = 24'b001011000010111000111001;
rgb[10276] = 24'b001110100011111001001101;
rgb[10277] = 24'b010010010100110101100000;
rgb[10278] = 24'b010110000101110101110011;
rgb[10279] = 24'b011001110110110110000110;
rgb[10280] = 24'b011110000111111010010111;
rgb[10281] = 24'b100010111001000010100110;
rgb[10282] = 24'b100111101010001010110101;
rgb[10283] = 24'b101100011011010111000100;
rgb[10284] = 24'b110001011100011111010010;
rgb[10285] = 24'b110110001101101011100001;
rgb[10286] = 24'b111010111110110011110000;
rgb[10287] = 24'b111111111111111111111111;
rgb[10288] = 24'b000000000000000000000000;
rgb[10289] = 24'b000011010000111000010100;
rgb[10290] = 24'b000110110001110100101000;
rgb[10291] = 24'b001010000010110000111101;
rgb[10292] = 24'b001101100011101101010001;
rgb[10293] = 24'b010001000100101001100101;
rgb[10294] = 24'b010100010101100101111010;
rgb[10295] = 24'b010111110110100010001110;
rgb[10296] = 24'b011100000111100110011111;
rgb[10297] = 24'b100001001000110010101101;
rgb[10298] = 24'b100110001001111110111011;
rgb[10299] = 24'b101011011011001011001000;
rgb[10300] = 24'b110000011100010111010110;
rgb[10301] = 24'b110101101101100011100011;
rgb[10302] = 24'b111010101110101111110001;
rgb[10303] = 24'b111111111111111111111111;
rgb[10304] = 24'b000000000000000000000000;
rgb[10305] = 24'b000011000000111000010101;
rgb[10306] = 24'b000110000001110000101011;
rgb[10307] = 24'b001001010010101001000000;
rgb[10308] = 24'b001100010011100001010110;
rgb[10309] = 24'b001111100100011001101011;
rgb[10310] = 24'b010010100101010110000001;
rgb[10311] = 24'b010101110110001110010110;
rgb[10312] = 24'b011010000111010010100111;
rgb[10313] = 24'b011111011000100010110100;
rgb[10314] = 24'b100100111001101111000000;
rgb[10315] = 24'b101010001010111111001101;
rgb[10316] = 24'b101111101100001111011001;
rgb[10317] = 24'b110100111101011111100110;
rgb[10318] = 24'b111010011110101111110010;
rgb[10319] = 24'b111111111111111111111111;
rgb[10320] = 24'b000000000000000000000000;
rgb[10321] = 24'b000010110000110100010110;
rgb[10322] = 24'b000101100001101000101101;
rgb[10323] = 24'b001000100010100001000100;
rgb[10324] = 24'b001011010011010101011010;
rgb[10325] = 24'b001110000100001101110001;
rgb[10326] = 24'b010001000101000010001000;
rgb[10327] = 24'b010011110101111010011110;
rgb[10328] = 24'b011000000110111110101111;
rgb[10329] = 24'b011101101000001110111011;
rgb[10330] = 24'b100011011001100011000110;
rgb[10331] = 24'b101001001010110011010001;
rgb[10332] = 24'b101110111100000111011101;
rgb[10333] = 24'b110100011101010111101000;
rgb[10334] = 24'b111010001110101011110011;
rgb[10335] = 24'b111111111111111111111111;
rgb[10336] = 24'b000000000000000000000000;
rgb[10337] = 24'b000010100000110000010111;
rgb[10338] = 24'b000101000001100100101111;
rgb[10339] = 24'b000111100010011001000111;
rgb[10340] = 24'b001010000011001101011111;
rgb[10341] = 24'b001100110011111101110110;
rgb[10342] = 24'b001111010100110010001110;
rgb[10343] = 24'b010001110101100110100110;
rgb[10344] = 24'b010110000110101010110111;
rgb[10345] = 24'b011100000111111111000001;
rgb[10346] = 24'b100001111001010011001100;
rgb[10347] = 24'b100111111010101011010110;
rgb[10348] = 24'b101101111011111111100000;
rgb[10349] = 24'b110011111101010011101010;
rgb[10350] = 24'b111001111110100111110100;
rgb[10351] = 24'b111111111111111111111110;
rgb[10352] = 24'b000000000000000000000000;
rgb[10353] = 24'b000010010000110000011000;
rgb[10354] = 24'b000100100001100000110001;
rgb[10355] = 24'b000110110010010001001010;
rgb[10356] = 24'b001001000011000001100011;
rgb[10357] = 24'b001011010011110001111100;
rgb[10358] = 24'b001101100100100010010101;
rgb[10359] = 24'b001111110101010010101110;
rgb[10360] = 24'b010100000110010110111111;
rgb[10361] = 24'b011010010111101111001000;
rgb[10362] = 24'b100000101001000111010001;
rgb[10363] = 24'b100110111010011111011010;
rgb[10364] = 24'b101101001011110111100011;
rgb[10365] = 24'b110011011101001111101100;
rgb[10366] = 24'b111001101110100111110101;
rgb[10367] = 24'b111111111111111111111111;
rgb[10368] = 24'b000000000000000000000000;
rgb[10369] = 24'b000001110000101100011010;
rgb[10370] = 24'b000011110001011000110100;
rgb[10371] = 24'b000101110010001001001110;
rgb[10372] = 24'b000111110010110101101000;
rgb[10373] = 24'b001001110011100010000010;
rgb[10374] = 24'b001011110100010010011100;
rgb[10375] = 24'b001101110100111110110110;
rgb[10376] = 24'b010010000110000011000111;
rgb[10377] = 24'b011000100111011111001111;
rgb[10378] = 24'b011111001000110111010111;
rgb[10379] = 24'b100101101010010011011111;
rgb[10380] = 24'b101100001011101111100111;
rgb[10381] = 24'b110010101101000111101111;
rgb[10382] = 24'b111001001110100011110111;
rgb[10383] = 24'b111111111111111111111110;
rgb[10384] = 24'b000000000000000000000000;
rgb[10385] = 24'b000001100000101000011011;
rgb[10386] = 24'b000011010001010100110110;
rgb[10387] = 24'b000101000010000001010001;
rgb[10388] = 24'b000110110010101001101100;
rgb[10389] = 24'b001000010011010110001000;
rgb[10390] = 24'b001010000100000010100011;
rgb[10391] = 24'b001011110100101010111110;
rgb[10392] = 24'b010000000101101111001111;
rgb[10393] = 24'b010110110111001111010110;
rgb[10394] = 24'b011101101000101011011101;
rgb[10395] = 24'b100100101010000111100011;
rgb[10396] = 24'b101011011011100111101010;
rgb[10397] = 24'b110010001101000011110001;
rgb[10398] = 24'b111000111110011111111000;
rgb[10399] = 24'b111111111111111111111111;
rgb[10400] = 24'b000000000000000000000000;
rgb[10401] = 24'b000001010000100100011100;
rgb[10402] = 24'b000010110001001100111000;
rgb[10403] = 24'b000100010001110101010101;
rgb[10404] = 24'b000101100010011101110001;
rgb[10405] = 24'b000111000011000110001101;
rgb[10406] = 24'b001000100011101110101010;
rgb[10407] = 24'b001001110100010111000110;
rgb[10408] = 24'b001110000101011011010111;
rgb[10409] = 24'b010101000110111011011101;
rgb[10410] = 24'b011100011000011011100010;
rgb[10411] = 24'b100011011001111011101000;
rgb[10412] = 24'b101010101011011011101110;
rgb[10413] = 24'b110001101100111011110011;
rgb[10414] = 24'b111000101110011011111001;
rgb[10415] = 24'b111111111111111111111110;
rgb[10416] = 24'b000000000000000000000000;
rgb[10417] = 24'b000001000000100100011101;
rgb[10418] = 24'b000010010001001000111010;
rgb[10419] = 24'b000011010001101101011000;
rgb[10420] = 24'b000100100010010101110101;
rgb[10421] = 24'b000101100010111010010011;
rgb[10422] = 24'b000110110011011110110000;
rgb[10423] = 24'b000111110100000011001110;
rgb[10424] = 24'b001100000101000111011111;
rgb[10425] = 24'b010011100110101011100011;
rgb[10426] = 24'b011010111000001111101000;
rgb[10427] = 24'b100010011001110011101100;
rgb[10428] = 24'b101001101011010011110001;
rgb[10429] = 24'b110001001100110111110101;
rgb[10430] = 24'b111000011110011011111010;
rgb[10431] = 24'b111111111111111111111111;
rgb[10432] = 24'b000000000000000000000000;
rgb[10433] = 24'b000000110000100000011110;
rgb[10434] = 24'b000001100001000100111101;
rgb[10435] = 24'b000010100001100101011011;
rgb[10436] = 24'b000011010010001001111010;
rgb[10437] = 24'b000100000010101010011001;
rgb[10438] = 24'b000101000011001110110111;
rgb[10439] = 24'b000101110011110011010110;
rgb[10440] = 24'b001010000100110111100111;
rgb[10441] = 24'b010001110110011011101010;
rgb[10442] = 24'b011001010111111111101110;
rgb[10443] = 24'b100001001001100111110001;
rgb[10444] = 24'b101000111011001011110100;
rgb[10445] = 24'b110000011100110011111000;
rgb[10446] = 24'b111000001110010111111011;
rgb[10447] = 24'b111111111111111111111111;
rgb[10448] = 24'b000000000000000000000000;
rgb[10449] = 24'b000000100000011100011111;
rgb[10450] = 24'b000001000000111100111111;
rgb[10451] = 24'b000001100001011101011111;
rgb[10452] = 24'b000010010001111101111110;
rgb[10453] = 24'b000010110010011110011110;
rgb[10454] = 24'b000011010010111110111110;
rgb[10455] = 24'b000011110011011111011110;
rgb[10456] = 24'b001000000100100011101111;
rgb[10457] = 24'b010000000110001011110001;
rgb[10458] = 24'b011000000111110011110011;
rgb[10459] = 24'b100000001001011011110101;
rgb[10460] = 24'b100111111011000011111000;
rgb[10461] = 24'b101111111100101011111010;
rgb[10462] = 24'b110111111110010011111100;
rgb[10463] = 24'b111111111111111111111111;
rgb[10464] = 24'b000000000000000000000000;
rgb[10465] = 24'b000000010000011100100000;
rgb[10466] = 24'b000000100000111001000001;
rgb[10467] = 24'b000000110001010101100010;
rgb[10468] = 24'b000001000001110010000011;
rgb[10469] = 24'b000001010010001110100100;
rgb[10470] = 24'b000001100010101111000101;
rgb[10471] = 24'b000001110011001011100110;
rgb[10472] = 24'b000110000100001111110111;
rgb[10473] = 24'b001110010101111011111000;
rgb[10474] = 24'b010110100111100011111001;
rgb[10475] = 24'b011110111001001111111010;
rgb[10476] = 24'b100111001010111011111011;
rgb[10477] = 24'b101111011100100111111100;
rgb[10478] = 24'b110111101110010011111101;
rgb[10479] = 24'b111111111111111111111111;
rgb[10480] = 24'b000000000000000000000000;
rgb[10481] = 24'b000000000000011000100010;
rgb[10482] = 24'b000000000000110001000100;
rgb[10483] = 24'b000000000001001101100110;
rgb[10484] = 24'b000000000001100110001000;
rgb[10485] = 24'b000000000010000010101010;
rgb[10486] = 24'b000000000010011011001100;
rgb[10487] = 24'b000000000010110111101110;
rgb[10488] = 24'b000100010011111011111110;
rgb[10489] = 24'b001100100101100111111111;
rgb[10490] = 24'b010101010111010111111110;
rgb[10491] = 24'b011101101001000011111111;
rgb[10492] = 24'b100110011010110011111111;
rgb[10493] = 24'b101110111100011111111111;
rgb[10494] = 24'b110111011110001111111111;
rgb[10495] = 24'b111111111111111111111111;
rgb[10496] = 24'b000000000000000000000000;
rgb[10497] = 24'b000100010001000100010001;
rgb[10498] = 24'b001000100010001000100010;
rgb[10499] = 24'b001100110011001100110011;
rgb[10500] = 24'b010001000100010001000100;
rgb[10501] = 24'b010101010101010101010101;
rgb[10502] = 24'b011001100110011001100110;
rgb[10503] = 24'b011101110111011101110111;
rgb[10504] = 24'b100010001000100010001000;
rgb[10505] = 24'b100110011001100110011001;
rgb[10506] = 24'b101010101010101010101010;
rgb[10507] = 24'b101110111011101110111011;
rgb[10508] = 24'b110011001100110011001100;
rgb[10509] = 24'b110111011101110111011101;
rgb[10510] = 24'b111011101110111011101110;
rgb[10511] = 24'b111111111111111111111111;
rgb[10512] = 24'b000000000000000000000000;
rgb[10513] = 24'b000011110001000000010010;
rgb[10514] = 24'b000111110010000000100100;
rgb[10515] = 24'b001011110011000000110110;
rgb[10516] = 24'b001111110100000001001000;
rgb[10517] = 24'b010011110101000001011010;
rgb[10518] = 24'b010111110110000001101100;
rgb[10519] = 24'b011011110111000001111110;
rgb[10520] = 24'b100000001000000110001111;
rgb[10521] = 24'b100100101001001110011111;
rgb[10522] = 24'b101001001010010110101111;
rgb[10523] = 24'b101101101011011110111111;
rgb[10524] = 24'b110010001100100111001111;
rgb[10525] = 24'b110110101101101111011111;
rgb[10526] = 24'b111011001110110111101111;
rgb[10527] = 24'b111111111111111111111111;
rgb[10528] = 24'b000000000000000000000000;
rgb[10529] = 24'b000011100000111100010011;
rgb[10530] = 24'b000111010001111000100110;
rgb[10531] = 24'b001011000010110100111001;
rgb[10532] = 24'b001110100011110001001101;
rgb[10533] = 24'b010010010100101101100000;
rgb[10534] = 24'b010110000101101001110011;
rgb[10535] = 24'b011001110110101010000110;
rgb[10536] = 24'b011110000111101110010111;
rgb[10537] = 24'b100010111000110110100110;
rgb[10538] = 24'b100111101010000010110101;
rgb[10539] = 24'b101100011011001111000100;
rgb[10540] = 24'b110001011100011011010010;
rgb[10541] = 24'b110110001101100111100001;
rgb[10542] = 24'b111010111110110011110000;
rgb[10543] = 24'b111111111111111111111111;
rgb[10544] = 24'b000000000000000000000000;
rgb[10545] = 24'b000011010000111000010100;
rgb[10546] = 24'b000110110001110000101000;
rgb[10547] = 24'b001010000010101000111101;
rgb[10548] = 24'b001101100011100001010001;
rgb[10549] = 24'b010001000100011101100101;
rgb[10550] = 24'b010100010101010101111010;
rgb[10551] = 24'b010111110110001110001110;
rgb[10552] = 24'b011100000111010010011111;
rgb[10553] = 24'b100001001000100010101101;
rgb[10554] = 24'b100110001001110010111011;
rgb[10555] = 24'b101011011010111111001000;
rgb[10556] = 24'b110000011100001111010110;
rgb[10557] = 24'b110101101101011111100011;
rgb[10558] = 24'b111010101110101111110001;
rgb[10559] = 24'b111111111111111111111111;
rgb[10560] = 24'b000000000000000000000000;
rgb[10561] = 24'b000011000000110100010101;
rgb[10562] = 24'b000110000001101000101011;
rgb[10563] = 24'b001001010010011101000000;
rgb[10564] = 24'b001100010011010101010110;
rgb[10565] = 24'b001111100100001001101011;
rgb[10566] = 24'b010010100100111110000001;
rgb[10567] = 24'b010101110101110110010110;
rgb[10568] = 24'b011010000110111010100111;
rgb[10569] = 24'b011111011000001010110100;
rgb[10570] = 24'b100100111001011111000000;
rgb[10571] = 24'b101010001010110011001101;
rgb[10572] = 24'b101111101100000011011001;
rgb[10573] = 24'b110100111101010111100110;
rgb[10574] = 24'b111010011110101011110010;
rgb[10575] = 24'b111111111111111111111111;
rgb[10576] = 24'b000000000000000000000000;
rgb[10577] = 24'b000010110000110000010110;
rgb[10578] = 24'b000101100001100000101101;
rgb[10579] = 24'b001000100010010101000100;
rgb[10580] = 24'b001011010011000101011010;
rgb[10581] = 24'b001110000011111001110001;
rgb[10582] = 24'b010001000100101010001000;
rgb[10583] = 24'b010011110101011010011110;
rgb[10584] = 24'b011000000110011110101111;
rgb[10585] = 24'b011101100111110110111011;
rgb[10586] = 24'b100011011001001111000110;
rgb[10587] = 24'b101001001010100011010001;
rgb[10588] = 24'b101110111011111011011101;
rgb[10589] = 24'b110100011101001111101000;
rgb[10590] = 24'b111010001110100111110011;
rgb[10591] = 24'b111111111111111111111111;
rgb[10592] = 24'b000000000000000000000000;
rgb[10593] = 24'b000010100000101100010111;
rgb[10594] = 24'b000101000001011000101111;
rgb[10595] = 24'b000111100010001001000111;
rgb[10596] = 24'b001010000010110101011111;
rgb[10597] = 24'b001100110011100101110110;
rgb[10598] = 24'b001111010100010010001110;
rgb[10599] = 24'b010001110101000010100110;
rgb[10600] = 24'b010110000110000110110111;
rgb[10601] = 24'b011100000111011111000001;
rgb[10602] = 24'b100001111000111011001100;
rgb[10603] = 24'b100111111010010011010110;
rgb[10604] = 24'b101101111011101111100000;
rgb[10605] = 24'b110011111101000111101010;
rgb[10606] = 24'b111001111110100011110100;
rgb[10607] = 24'b111111111111111111111110;
rgb[10608] = 24'b000000000000000000000000;
rgb[10609] = 24'b000010010000101000011000;
rgb[10610] = 24'b000100100001010100110001;
rgb[10611] = 24'b000110110001111101001010;
rgb[10612] = 24'b001001000010101001100011;
rgb[10613] = 24'b001011010011010001111100;
rgb[10614] = 24'b001101100011111110010101;
rgb[10615] = 24'b001111110100101010101110;
rgb[10616] = 24'b010100000101101110111111;
rgb[10617] = 24'b011010010111001011001000;
rgb[10618] = 24'b100000101000100111010001;
rgb[10619] = 24'b100110111010000111011010;
rgb[10620] = 24'b101101001011100011100011;
rgb[10621] = 24'b110011011101000011101100;
rgb[10622] = 24'b111001101110011111110101;
rgb[10623] = 24'b111111111111111111111111;
rgb[10624] = 24'b000000000000000000000000;
rgb[10625] = 24'b000001110000100100011010;
rgb[10626] = 24'b000011110001001100110100;
rgb[10627] = 24'b000101110001110001001110;
rgb[10628] = 24'b000111110010011001101000;
rgb[10629] = 24'b001001110011000010000010;
rgb[10630] = 24'b001011110011100110011100;
rgb[10631] = 24'b001101110100001110110110;
rgb[10632] = 24'b010010000101010011000111;
rgb[10633] = 24'b011000100110110011001111;
rgb[10634] = 24'b011111001000010111010111;
rgb[10635] = 24'b100101101001110111011111;
rgb[10636] = 24'b101100001011010111100111;
rgb[10637] = 24'b110010101100111011101111;
rgb[10638] = 24'b111001001110011011110111;
rgb[10639] = 24'b111111111111111111111110;
rgb[10640] = 24'b000000000000000000000000;
rgb[10641] = 24'b000001100000100000011011;
rgb[10642] = 24'b000011010001000100110110;
rgb[10643] = 24'b000101000001101001010001;
rgb[10644] = 24'b000110110010001001101100;
rgb[10645] = 24'b001000010010101110001000;
rgb[10646] = 24'b001010000011010010100011;
rgb[10647] = 24'b001011110011110110111110;
rgb[10648] = 24'b010000000100111011001111;
rgb[10649] = 24'b010110110110011111010110;
rgb[10650] = 24'b011101101000000011011101;
rgb[10651] = 24'b100100101001100111100011;
rgb[10652] = 24'b101011011011001111101010;
rgb[10653] = 24'b110010001100110011110001;
rgb[10654] = 24'b111000111110010111111000;
rgb[10655] = 24'b111111111111111111111111;
rgb[10656] = 24'b000000000000000000000000;
rgb[10657] = 24'b000001010000011100011100;
rgb[10658] = 24'b000010110000111100111000;
rgb[10659] = 24'b000100010001011101010101;
rgb[10660] = 24'b000101100001111101110001;
rgb[10661] = 24'b000111000010011110001101;
rgb[10662] = 24'b001000100010111010101010;
rgb[10663] = 24'b001001110011011011000110;
rgb[10664] = 24'b001110000100011111010111;
rgb[10665] = 24'b010101000110000111011101;
rgb[10666] = 24'b011100010111110011100010;
rgb[10667] = 24'b100011011001011011101000;
rgb[10668] = 24'b101010101011000011101110;
rgb[10669] = 24'b110001101100101011110011;
rgb[10670] = 24'b111000101110010011111001;
rgb[10671] = 24'b111111111111111111111110;
rgb[10672] = 24'b000000000000000000000000;
rgb[10673] = 24'b000001000000011000011101;
rgb[10674] = 24'b000010010000110100111010;
rgb[10675] = 24'b000011010001010001011000;
rgb[10676] = 24'b000100100001101101110101;
rgb[10677] = 24'b000101100010001010010011;
rgb[10678] = 24'b000110110010100110110000;
rgb[10679] = 24'b000111110011000011001110;
rgb[10680] = 24'b001100000100000111011111;
rgb[10681] = 24'b010011100101110011100011;
rgb[10682] = 24'b011010110111011111101000;
rgb[10683] = 24'b100010011001001011101100;
rgb[10684] = 24'b101001101010110111110001;
rgb[10685] = 24'b110001001100100011110101;
rgb[10686] = 24'b111000011110001111111010;
rgb[10687] = 24'b111111111111111111111111;
rgb[10688] = 24'b000000000000000000000000;
rgb[10689] = 24'b000000110000010100011110;
rgb[10690] = 24'b000001100000101100111101;
rgb[10691] = 24'b000010100001000101011011;
rgb[10692] = 24'b000011010001011101111010;
rgb[10693] = 24'b000100000001110110011001;
rgb[10694] = 24'b000101000010001110110111;
rgb[10695] = 24'b000101110010100111010110;
rgb[10696] = 24'b001010000011101011100111;
rgb[10697] = 24'b010001110101011011101010;
rgb[10698] = 24'b011001010111001011101110;
rgb[10699] = 24'b100001001000111011110001;
rgb[10700] = 24'b101000111010101011110100;
rgb[10701] = 24'b110000011100011011111000;
rgb[10702] = 24'b111000001110001011111011;
rgb[10703] = 24'b111111111111111111111111;
rgb[10704] = 24'b000000000000000000000000;
rgb[10705] = 24'b000000100000010100011111;
rgb[10706] = 24'b000001000000101000111111;
rgb[10707] = 24'b000001100000111101011111;
rgb[10708] = 24'b000010010001010001111110;
rgb[10709] = 24'b000010110001100110011110;
rgb[10710] = 24'b000011010001111010111110;
rgb[10711] = 24'b000011110010001111011110;
rgb[10712] = 24'b001000000011010011101111;
rgb[10713] = 24'b010000000101000111110001;
rgb[10714] = 24'b011000000110111011110011;
rgb[10715] = 24'b100000001000101111110101;
rgb[10716] = 24'b100111111010100011111000;
rgb[10717] = 24'b101111111100010111111010;
rgb[10718] = 24'b110111111110001011111100;
rgb[10719] = 24'b111111111111111111111111;
rgb[10720] = 24'b000000000000000000000000;
rgb[10721] = 24'b000000010000010000100000;
rgb[10722] = 24'b000000100000100001000001;
rgb[10723] = 24'b000000110000110001100010;
rgb[10724] = 24'b000001000001000010000011;
rgb[10725] = 24'b000001010001010010100100;
rgb[10726] = 24'b000001100001100011000101;
rgb[10727] = 24'b000001110001110111100110;
rgb[10728] = 24'b000110000010111011110111;
rgb[10729] = 24'b001110010100101111111000;
rgb[10730] = 24'b010110100110100111111001;
rgb[10731] = 24'b011110111000011111111010;
rgb[10732] = 24'b100111001010010111111011;
rgb[10733] = 24'b101111011100001111111100;
rgb[10734] = 24'b110111101110000111111101;
rgb[10735] = 24'b111111111111111111111111;
rgb[10736] = 24'b000000000000000000000000;
rgb[10737] = 24'b000000000000001100100010;
rgb[10738] = 24'b000000000000011001000100;
rgb[10739] = 24'b000000000000100101100110;
rgb[10740] = 24'b000000000000110010001000;
rgb[10741] = 24'b000000000001000010101010;
rgb[10742] = 24'b000000000001001111001100;
rgb[10743] = 24'b000000000001011011101110;
rgb[10744] = 24'b000100010010011111111110;
rgb[10745] = 24'b001100100100011011111111;
rgb[10746] = 24'b010101010110010111111110;
rgb[10747] = 24'b011101101000001111111111;
rgb[10748] = 24'b100110011010001011111111;
rgb[10749] = 24'b101110111100000111111111;
rgb[10750] = 24'b110111011110000011111111;
rgb[10751] = 24'b111111111111111111111111;
rgb[10752] = 24'b000000000000000000000000;
rgb[10753] = 24'b000100010001000100010001;
rgb[10754] = 24'b001000100010001000100010;
rgb[10755] = 24'b001100110011001100110011;
rgb[10756] = 24'b010001000100010001000100;
rgb[10757] = 24'b010101010101010101010101;
rgb[10758] = 24'b011001100110011001100110;
rgb[10759] = 24'b011101110111011101110111;
rgb[10760] = 24'b100010001000100010001000;
rgb[10761] = 24'b100110011001100110011001;
rgb[10762] = 24'b101010101010101010101010;
rgb[10763] = 24'b101110111011101110111011;
rgb[10764] = 24'b110011001100110011001100;
rgb[10765] = 24'b110111011101110111011101;
rgb[10766] = 24'b111011101110111011101110;
rgb[10767] = 24'b111111111111111111111111;
rgb[10768] = 24'b000000000000000000000000;
rgb[10769] = 24'b000011110000111100010010;
rgb[10770] = 24'b000111110001111100100100;
rgb[10771] = 24'b001011110010111100110110;
rgb[10772] = 24'b001111110011111101001000;
rgb[10773] = 24'b010011110100111101011010;
rgb[10774] = 24'b010111110101111101101100;
rgb[10775] = 24'b011011110110111101111110;
rgb[10776] = 24'b100000001000000010001111;
rgb[10777] = 24'b100100101001001010011111;
rgb[10778] = 24'b101001001010010010101111;
rgb[10779] = 24'b101101101011011010111111;
rgb[10780] = 24'b110010001100100011001111;
rgb[10781] = 24'b110110101101101011011111;
rgb[10782] = 24'b111011001110110011101111;
rgb[10783] = 24'b111111111111111111111111;
rgb[10784] = 24'b000000000000000000000000;
rgb[10785] = 24'b000011100000111000010011;
rgb[10786] = 24'b000111010001110100100110;
rgb[10787] = 24'b001011000010110000111001;
rgb[10788] = 24'b001110100011101001001101;
rgb[10789] = 24'b010010010100100101100000;
rgb[10790] = 24'b010110000101100001110011;
rgb[10791] = 24'b011001110110011110000110;
rgb[10792] = 24'b011110000111100010010111;
rgb[10793] = 24'b100010111000101110100110;
rgb[10794] = 24'b100111101001111010110101;
rgb[10795] = 24'b101100011011000111000100;
rgb[10796] = 24'b110001011100010111010010;
rgb[10797] = 24'b110110001101100011100001;
rgb[10798] = 24'b111010111110101111110000;
rgb[10799] = 24'b111111111111111111111111;
rgb[10800] = 24'b000000000000000000000000;
rgb[10801] = 24'b000011010000110100010100;
rgb[10802] = 24'b000110110001101100101000;
rgb[10803] = 24'b001010000010100000111101;
rgb[10804] = 24'b001101100011011001010001;
rgb[10805] = 24'b010001000100010001100101;
rgb[10806] = 24'b010100010101000101111010;
rgb[10807] = 24'b010111110101111110001110;
rgb[10808] = 24'b011100000111000010011111;
rgb[10809] = 24'b100001001000010010101101;
rgb[10810] = 24'b100110001001100010111011;
rgb[10811] = 24'b101011011010110111001000;
rgb[10812] = 24'b110000011100000111010110;
rgb[10813] = 24'b110101101101011011100011;
rgb[10814] = 24'b111010101110101011110001;
rgb[10815] = 24'b111111111111111111111111;
rgb[10816] = 24'b000000000000000000000000;
rgb[10817] = 24'b000011000000110000010101;
rgb[10818] = 24'b000110000001100000101011;
rgb[10819] = 24'b001001010010010101000000;
rgb[10820] = 24'b001100010011000101010110;
rgb[10821] = 24'b001111100011111001101011;
rgb[10822] = 24'b010010100100101010000001;
rgb[10823] = 24'b010101110101011110010110;
rgb[10824] = 24'b011010000110100010100111;
rgb[10825] = 24'b011111010111110110110100;
rgb[10826] = 24'b100100111001001111000000;
rgb[10827] = 24'b101010001010100011001101;
rgb[10828] = 24'b101111101011111011011001;
rgb[10829] = 24'b110100111101001111100110;
rgb[10830] = 24'b111010011110100111110010;
rgb[10831] = 24'b111111111111111111111111;
rgb[10832] = 24'b000000000000000000000000;
rgb[10833] = 24'b000010110000101100010110;
rgb[10834] = 24'b000101100001011000101101;
rgb[10835] = 24'b001000100010001001000100;
rgb[10836] = 24'b001011010010110101011010;
rgb[10837] = 24'b001110000011100001110001;
rgb[10838] = 24'b010001000100010010001000;
rgb[10839] = 24'b010011110100111110011110;
rgb[10840] = 24'b011000000110000010101111;
rgb[10841] = 24'b011101100111011010111011;
rgb[10842] = 24'b100011011000110111000110;
rgb[10843] = 24'b101001001010010011010001;
rgb[10844] = 24'b101110111011101111011101;
rgb[10845] = 24'b110100011101000111101000;
rgb[10846] = 24'b111010001110100011110011;
rgb[10847] = 24'b111111111111111111111111;
rgb[10848] = 24'b000000000000000000000000;
rgb[10849] = 24'b000010100000101000010111;
rgb[10850] = 24'b000101000001010000101111;
rgb[10851] = 24'b000111100001111001000111;
rgb[10852] = 24'b001010000010100001011111;
rgb[10853] = 24'b001100110011001101110110;
rgb[10854] = 24'b001111010011110110001110;
rgb[10855] = 24'b010001110100011110100110;
rgb[10856] = 24'b010110000101100010110111;
rgb[10857] = 24'b011100000111000011000001;
rgb[10858] = 24'b100001111000011111001100;
rgb[10859] = 24'b100111111001111111010110;
rgb[10860] = 24'b101101111011011111100000;
rgb[10861] = 24'b110011111100111111101010;
rgb[10862] = 24'b111001111110011111110100;
rgb[10863] = 24'b111111111111111111111110;
rgb[10864] = 24'b000000000000000000000000;
rgb[10865] = 24'b000010010000100100011000;
rgb[10866] = 24'b000100100001001000110001;
rgb[10867] = 24'b000110110001101101001010;
rgb[10868] = 24'b001001000010010001100011;
rgb[10869] = 24'b001011010010110101111100;
rgb[10870] = 24'b001101100011011010010101;
rgb[10871] = 24'b001111110011111110101110;
rgb[10872] = 24'b010100000101000010111111;
rgb[10873] = 24'b011010010110100111001000;
rgb[10874] = 24'b100000101000001011010001;
rgb[10875] = 24'b100110111001101111011010;
rgb[10876] = 24'b101101001011010011100011;
rgb[10877] = 24'b110011011100110111101100;
rgb[10878] = 24'b111001101110011011110101;
rgb[10879] = 24'b111111111111111111111111;
rgb[10880] = 24'b000000000000000000000000;
rgb[10881] = 24'b000001110000011100011010;
rgb[10882] = 24'b000011110000111100110100;
rgb[10883] = 24'b000101110001011101001110;
rgb[10884] = 24'b000111110001111101101000;
rgb[10885] = 24'b001001110010011110000010;
rgb[10886] = 24'b001011110010111110011100;
rgb[10887] = 24'b001101110011011110110110;
rgb[10888] = 24'b010010000100100011000111;
rgb[10889] = 24'b011000100110001011001111;
rgb[10890] = 24'b011111000111110011010111;
rgb[10891] = 24'b100101101001011011011111;
rgb[10892] = 24'b101100001011000011100111;
rgb[10893] = 24'b110010101100101011101111;
rgb[10894] = 24'b111001001110010011110111;
rgb[10895] = 24'b111111111111111111111110;
rgb[10896] = 24'b000000000000000000000000;
rgb[10897] = 24'b000001100000011000011011;
rgb[10898] = 24'b000011010000110100110110;
rgb[10899] = 24'b000101000001010001010001;
rgb[10900] = 24'b000110110001101101101100;
rgb[10901] = 24'b001000010010000110001000;
rgb[10902] = 24'b001010000010100010100011;
rgb[10903] = 24'b001011110010111110111110;
rgb[10904] = 24'b010000000100000011001111;
rgb[10905] = 24'b010110110101101111010110;
rgb[10906] = 24'b011101100111011011011101;
rgb[10907] = 24'b100100101001001011100011;
rgb[10908] = 24'b101011011010110111101010;
rgb[10909] = 24'b110010001100100011110001;
rgb[10910] = 24'b111000111110001111111000;
rgb[10911] = 24'b111111111111111111111111;
rgb[10912] = 24'b000000000000000000000000;
rgb[10913] = 24'b000001010000010100011100;
rgb[10914] = 24'b000010110000101100111000;
rgb[10915] = 24'b000100010001000101010101;
rgb[10916] = 24'b000101100001011001110001;
rgb[10917] = 24'b000111000001110010001101;
rgb[10918] = 24'b001000100010001010101010;
rgb[10919] = 24'b001001110010011111000110;
rgb[10920] = 24'b001110000011100011010111;
rgb[10921] = 24'b010101000101010011011101;
rgb[10922] = 24'b011100010111000111100010;
rgb[10923] = 24'b100011011000110111101000;
rgb[10924] = 24'b101010101010101011101110;
rgb[10925] = 24'b110001101100011011110011;
rgb[10926] = 24'b111000101110001011111001;
rgb[10927] = 24'b111111111111111111111110;
rgb[10928] = 24'b000000000000000000000000;
rgb[10929] = 24'b000001000000010000011101;
rgb[10930] = 24'b000010010000100100111010;
rgb[10931] = 24'b000011010000110101011000;
rgb[10932] = 24'b000100100001001001110101;
rgb[10933] = 24'b000101100001011010010011;
rgb[10934] = 24'b000110110001101110110000;
rgb[10935] = 24'b000111110001111111001110;
rgb[10936] = 24'b001100000011000011011111;
rgb[10937] = 24'b010011100100111011100011;
rgb[10938] = 24'b011010110110101111101000;
rgb[10939] = 24'b100010011000100111101100;
rgb[10940] = 24'b101001101010011011110001;
rgb[10941] = 24'b110001001100010011110101;
rgb[10942] = 24'b111000011110000111111010;
rgb[10943] = 24'b111111111111111111111111;
rgb[10944] = 24'b000000000000000000000000;
rgb[10945] = 24'b000000110000001100011110;
rgb[10946] = 24'b000001100000011000111101;
rgb[10947] = 24'b000010100000101001011011;
rgb[10948] = 24'b000011010000110101111010;
rgb[10949] = 24'b000100000001000010011001;
rgb[10950] = 24'b000101000001010010110111;
rgb[10951] = 24'b000101110001011111010110;
rgb[10952] = 24'b001010000010100011100111;
rgb[10953] = 24'b010001110100011111101010;
rgb[10954] = 24'b011001010110010111101110;
rgb[10955] = 24'b100001001000010011110001;
rgb[10956] = 24'b101000111010001111110100;
rgb[10957] = 24'b110000011100000111111000;
rgb[10958] = 24'b111000001110000011111011;
rgb[10959] = 24'b111111111111111111111111;
rgb[10960] = 24'b000000000000000000000000;
rgb[10961] = 24'b000000100000001000011111;
rgb[10962] = 24'b000001000000010000111111;
rgb[10963] = 24'b000001100000011001011111;
rgb[10964] = 24'b000010010000100101111110;
rgb[10965] = 24'b000010110000101110011110;
rgb[10966] = 24'b000011010000110110111110;
rgb[10967] = 24'b000011110000111111011110;
rgb[10968] = 24'b001000000010000011101111;
rgb[10969] = 24'b010000000100000011110001;
rgb[10970] = 24'b011000000110000011110011;
rgb[10971] = 24'b100000001000000011110101;
rgb[10972] = 24'b100111111001111111111000;
rgb[10973] = 24'b101111111011111111111010;
rgb[10974] = 24'b110111111101111111111100;
rgb[10975] = 24'b111111111111111111111111;
rgb[10976] = 24'b000000000000000000000000;
rgb[10977] = 24'b000000010000000100100000;
rgb[10978] = 24'b000000100000001001000001;
rgb[10979] = 24'b000000110000001101100010;
rgb[10980] = 24'b000001000000010010000011;
rgb[10981] = 24'b000001010000010110100100;
rgb[10982] = 24'b000001100000011011000101;
rgb[10983] = 24'b000001110000011111100110;
rgb[10984] = 24'b000110000001100011110111;
rgb[10985] = 24'b001110010011100111111000;
rgb[10986] = 24'b010110100101101011111001;
rgb[10987] = 24'b011110110111101111111010;
rgb[10988] = 24'b100111001001110011111011;
rgb[10989] = 24'b101111011011110111111100;
rgb[10990] = 24'b110111101101111011111101;
rgb[10991] = 24'b111111111111111111111111;
rgb[10992] = 24'b000000000000000000000000;
rgb[10993] = 24'b000000000000000000100010;
rgb[10994] = 24'b000000000000000001000100;
rgb[10995] = 24'b000000000000000001100110;
rgb[10996] = 24'b000000000000000010001000;
rgb[10997] = 24'b000000000000000010101010;
rgb[10998] = 24'b000000000000000011001100;
rgb[10999] = 24'b000000000000000011101110;
rgb[11000] = 24'b000100010001000111111110;
rgb[11001] = 24'b001100100011001011111111;
rgb[11002] = 24'b010101010101010111111110;
rgb[11003] = 24'b011101100111011011111111;
rgb[11004] = 24'b100110011001100111111111;
rgb[11005] = 24'b101110111011101111111111;
rgb[11006] = 24'b110111011101110111111111;
rgb[11007] = 24'b111111111111111111111111;
rgb[11008] = 24'b000000000000000000000000;
rgb[11009] = 24'b000100010001000100010001;
rgb[11010] = 24'b001000100010001000100010;
rgb[11011] = 24'b001100110011001100110011;
rgb[11012] = 24'b010001000100010001000100;
rgb[11013] = 24'b010101010101010101010101;
rgb[11014] = 24'b011001100110011001100110;
rgb[11015] = 24'b011101110111011101110111;
rgb[11016] = 24'b100010001000100010001000;
rgb[11017] = 24'b100110011001100110011001;
rgb[11018] = 24'b101010101010101010101010;
rgb[11019] = 24'b101110111011101110111011;
rgb[11020] = 24'b110011001100110011001100;
rgb[11021] = 24'b110111011101110111011101;
rgb[11022] = 24'b111011101110111011101110;
rgb[11023] = 24'b111111111111111111111111;
rgb[11024] = 24'b000000000000000000000000;
rgb[11025] = 24'b000100000000111100010010;
rgb[11026] = 24'b001000000001111100100100;
rgb[11027] = 24'b001100000010111100110110;
rgb[11028] = 24'b010000000011111101001000;
rgb[11029] = 24'b010100000100111101011010;
rgb[11030] = 24'b011000000101111101101100;
rgb[11031] = 24'b011100000110111101111110;
rgb[11032] = 24'b100000011000000010001111;
rgb[11033] = 24'b100100111001001010011111;
rgb[11034] = 24'b101001011010010010101111;
rgb[11035] = 24'b101101111011011010111111;
rgb[11036] = 24'b110010011100100011001111;
rgb[11037] = 24'b110110111101101011011111;
rgb[11038] = 24'b111011011110110011101111;
rgb[11039] = 24'b111111111111111111111111;
rgb[11040] = 24'b000000000000000000000000;
rgb[11041] = 24'b000011110000111000010011;
rgb[11042] = 24'b000111100001110100100110;
rgb[11043] = 24'b001011010010110000111001;
rgb[11044] = 24'b001111000011101001001101;
rgb[11045] = 24'b010010110100100101100000;
rgb[11046] = 24'b010110100101100001110011;
rgb[11047] = 24'b011010100110011110000110;
rgb[11048] = 24'b011110110111100010010111;
rgb[11049] = 24'b100011011000101110100110;
rgb[11050] = 24'b101000001001111010110101;
rgb[11051] = 24'b101100111011000111000100;
rgb[11052] = 24'b110001101100010111010010;
rgb[11053] = 24'b110110011101100011100001;
rgb[11054] = 24'b111011001110101111110000;
rgb[11055] = 24'b111111111111111111111111;
rgb[11056] = 24'b000000000000000000000000;
rgb[11057] = 24'b000011100000110100010100;
rgb[11058] = 24'b000111000001101100101000;
rgb[11059] = 24'b001010100010100000111101;
rgb[11060] = 24'b001110000011011001010001;
rgb[11061] = 24'b010001110100010001100101;
rgb[11062] = 24'b010101010101000101111010;
rgb[11063] = 24'b011000110101111110001110;
rgb[11064] = 24'b011101000111000010011111;
rgb[11065] = 24'b100010001000010010101101;
rgb[11066] = 24'b100111001001100010111011;
rgb[11067] = 24'b101011111010110111001000;
rgb[11068] = 24'b110000111100000111010110;
rgb[11069] = 24'b110101111101011011100011;
rgb[11070] = 24'b111010111110101011110001;
rgb[11071] = 24'b111111111111111111111111;
rgb[11072] = 24'b000000000000000000000000;
rgb[11073] = 24'b000011010000110000010101;
rgb[11074] = 24'b000110100001100000101011;
rgb[11075] = 24'b001001110010010101000000;
rgb[11076] = 24'b001101010011000101010110;
rgb[11077] = 24'b010000100011111001101011;
rgb[11078] = 24'b010011110100101010000001;
rgb[11079] = 24'b010111010101011110010110;
rgb[11080] = 24'b011011100110100010100111;
rgb[11081] = 24'b100000100111110110110100;
rgb[11082] = 24'b100101111001001111000000;
rgb[11083] = 24'b101011001010100011001101;
rgb[11084] = 24'b110000001011111011011001;
rgb[11085] = 24'b110101011101001111100110;
rgb[11086] = 24'b111010101110100111110010;
rgb[11087] = 24'b111111111111111111111111;
rgb[11088] = 24'b000000000000000000000000;
rgb[11089] = 24'b000011000000101100010110;
rgb[11090] = 24'b000110000001011000101101;
rgb[11091] = 24'b001001010010001001000100;
rgb[11092] = 24'b001100010010110101011010;
rgb[11093] = 24'b001111100011100001110001;
rgb[11094] = 24'b010010100100010010001000;
rgb[11095] = 24'b010101100100111110011110;
rgb[11096] = 24'b011001110110000010101111;
rgb[11097] = 24'b011111010111011010111011;
rgb[11098] = 24'b100100111000110111000110;
rgb[11099] = 24'b101010001010010011010001;
rgb[11100] = 24'b101111101011101111011101;
rgb[11101] = 24'b110100111101000111101000;
rgb[11102] = 24'b111010011110100011110011;
rgb[11103] = 24'b111111111111111111111111;
rgb[11104] = 24'b000000000000000000000000;
rgb[11105] = 24'b000010110000101000010111;
rgb[11106] = 24'b000101100001010000101111;
rgb[11107] = 24'b001000100001111001000111;
rgb[11108] = 24'b001011010010100001011111;
rgb[11109] = 24'b001110010011001101110110;
rgb[11110] = 24'b010001000011110110001110;
rgb[11111] = 24'b010100000100011110100110;
rgb[11112] = 24'b011000010101100010110111;
rgb[11113] = 24'b011101110111000011000001;
rgb[11114] = 24'b100011101000011111001100;
rgb[11115] = 24'b101001001001111111010110;
rgb[11116] = 24'b101110111011011111100000;
rgb[11117] = 24'b110100011100111111101010;
rgb[11118] = 24'b111010001110011111110100;
rgb[11119] = 24'b111111111111111111111110;
rgb[11120] = 24'b000000000000000000000000;
rgb[11121] = 24'b000010100000100100011000;
rgb[11122] = 24'b000101010001001000110001;
rgb[11123] = 24'b000111110001101101001010;
rgb[11124] = 24'b001010100010010001100011;
rgb[11125] = 24'b001101000010110101111100;
rgb[11126] = 24'b001111110011011010010101;
rgb[11127] = 24'b010010100011111110101110;
rgb[11128] = 24'b010110110101000010111111;
rgb[11129] = 24'b011100100110100111001000;
rgb[11130] = 24'b100010011000001011010001;
rgb[11131] = 24'b101000011001101111011010;
rgb[11132] = 24'b101110001011010011100011;
rgb[11133] = 24'b110100001100110111101100;
rgb[11134] = 24'b111001111110011011110101;
rgb[11135] = 24'b111111111111111111111111;
rgb[11136] = 24'b000000000000000000000000;
rgb[11137] = 24'b000010010000011100011010;
rgb[11138] = 24'b000100110000111100110100;
rgb[11139] = 24'b000111000001011101001110;
rgb[11140] = 24'b001001100001111101101000;
rgb[11141] = 24'b001100000010011110000010;
rgb[11142] = 24'b001110010010111110011100;
rgb[11143] = 24'b010000110011011110110110;
rgb[11144] = 24'b010101000100100011000111;
rgb[11145] = 24'b011011000110001011001111;
rgb[11146] = 24'b100001010111110011010111;
rgb[11147] = 24'b100111011001011011011111;
rgb[11148] = 24'b101101011011000011100111;
rgb[11149] = 24'b110011101100101011101111;
rgb[11150] = 24'b111001101110010011110111;
rgb[11151] = 24'b111111111111111111111110;
rgb[11152] = 24'b000000000000000000000000;
rgb[11153] = 24'b000010000000011000011011;
rgb[11154] = 24'b000100010000110100110110;
rgb[11155] = 24'b000110100001010001010001;
rgb[11156] = 24'b001000100001101101101100;
rgb[11157] = 24'b001010110010000110001000;
rgb[11158] = 24'b001101000010100010100011;
rgb[11159] = 24'b001111010010111110111110;
rgb[11160] = 24'b010011100100000011001111;
rgb[11161] = 24'b011001110101101111010110;
rgb[11162] = 24'b100000000111011011011101;
rgb[11163] = 24'b100110011001001011100011;
rgb[11164] = 24'b101100111010110111101010;
rgb[11165] = 24'b110011001100100011110001;
rgb[11166] = 24'b111001011110001111111000;
rgb[11167] = 24'b111111111111111111111111;
rgb[11168] = 24'b000000000000000000000000;
rgb[11169] = 24'b000001110000010100011100;
rgb[11170] = 24'b000011110000101100111000;
rgb[11171] = 24'b000101110001000101010101;
rgb[11172] = 24'b000111110001011001110001;
rgb[11173] = 24'b001001110001110010001101;
rgb[11174] = 24'b001011100010001010101010;
rgb[11175] = 24'b001101100010011111000110;
rgb[11176] = 24'b010001110011100011010111;
rgb[11177] = 24'b011000010101010011011101;
rgb[11178] = 24'b011111000111000111100010;
rgb[11179] = 24'b100101101000110111101000;
rgb[11180] = 24'b101100001010101011101110;
rgb[11181] = 24'b110010101100011011110011;
rgb[11182] = 24'b111001001110001011111001;
rgb[11183] = 24'b111111111111111111111110;
rgb[11184] = 24'b000000000000000000000000;
rgb[11185] = 24'b000001100000010000011101;
rgb[11186] = 24'b000011010000100100111010;
rgb[11187] = 24'b000101000000110101011000;
rgb[11188] = 24'b000110110001001001110101;
rgb[11189] = 24'b001000100001011010010011;
rgb[11190] = 24'b001010010001101110110000;
rgb[11191] = 24'b001100000001111111001110;
rgb[11192] = 24'b010000010011000011011111;
rgb[11193] = 24'b010111000100111011100011;
rgb[11194] = 24'b011101110110101111101000;
rgb[11195] = 24'b100100101000100111101100;
rgb[11196] = 24'b101011011010011011110001;
rgb[11197] = 24'b110010001100010011110101;
rgb[11198] = 24'b111000111110000111111010;
rgb[11199] = 24'b111111111111111111111111;
rgb[11200] = 24'b000000000000000000000000;
rgb[11201] = 24'b000001010000001100011110;
rgb[11202] = 24'b000010110000011000111101;
rgb[11203] = 24'b000100010000101001011011;
rgb[11204] = 24'b000101110000110101111010;
rgb[11205] = 24'b000111010001000010011001;
rgb[11206] = 24'b001000110001010010110111;
rgb[11207] = 24'b001010010001011111010110;
rgb[11208] = 24'b001110100010100011100111;
rgb[11209] = 24'b010101100100011111101010;
rgb[11210] = 24'b011100100110010111101110;
rgb[11211] = 24'b100011101000010011110001;
rgb[11212] = 24'b101010101010001111110100;
rgb[11213] = 24'b110001101100000111111000;
rgb[11214] = 24'b111000101110000011111011;
rgb[11215] = 24'b111111111111111111111111;
rgb[11216] = 24'b000000000000000000000000;
rgb[11217] = 24'b000001010000001000011111;
rgb[11218] = 24'b000010100000010000111111;
rgb[11219] = 24'b000011110000011001011111;
rgb[11220] = 24'b000101000000100101111110;
rgb[11221] = 24'b000110010000101110011110;
rgb[11222] = 24'b000111100000110110111110;
rgb[11223] = 24'b001000110000111111011110;
rgb[11224] = 24'b001101000010000011101111;
rgb[11225] = 24'b010100010100000011110001;
rgb[11226] = 24'b011011100110000011110011;
rgb[11227] = 24'b100010111000000011110101;
rgb[11228] = 24'b101010001001111111111000;
rgb[11229] = 24'b110001011011111111111010;
rgb[11230] = 24'b111000101101111111111100;
rgb[11231] = 24'b111111111111111111111111;
rgb[11232] = 24'b000000000000000000000000;
rgb[11233] = 24'b000001000000000100100000;
rgb[11234] = 24'b000010000000001001000001;
rgb[11235] = 24'b000011000000001101100010;
rgb[11236] = 24'b000100000000010010000011;
rgb[11237] = 24'b000101000000010110100100;
rgb[11238] = 24'b000110000000011011000101;
rgb[11239] = 24'b000111010000011111100110;
rgb[11240] = 24'b001011100001100011110111;
rgb[11241] = 24'b010010110011100111111000;
rgb[11242] = 24'b011010010101101011111001;
rgb[11243] = 24'b100001110111101111111010;
rgb[11244] = 24'b101001011001110011111011;
rgb[11245] = 24'b110000111011110111111100;
rgb[11246] = 24'b111000011101111011111101;
rgb[11247] = 24'b111111111111111111111111;
rgb[11248] = 24'b000000000000000000000000;
rgb[11249] = 24'b000000110000000000100010;
rgb[11250] = 24'b000001100000000001000100;
rgb[11251] = 24'b000010010000000001100110;
rgb[11252] = 24'b000011000000000010001000;
rgb[11253] = 24'b000100000000000010101010;
rgb[11254] = 24'b000100110000000011001100;
rgb[11255] = 24'b000101100000000011101110;
rgb[11256] = 24'b001001110001000111111110;
rgb[11257] = 24'b010001100011001011111111;
rgb[11258] = 24'b011001010101010111111110;
rgb[11259] = 24'b100000110111011011111111;
rgb[11260] = 24'b101000101001100111111111;
rgb[11261] = 24'b110000011011101111111111;
rgb[11262] = 24'b111000001101110111111111;
rgb[11263] = 24'b111111111111111111111111;
rgb[11264] = 24'b000000000000000000000000;
rgb[11265] = 24'b000100010001000100010001;
rgb[11266] = 24'b001000100010001000100010;
rgb[11267] = 24'b001100110011001100110011;
rgb[11268] = 24'b010001000100010001000100;
rgb[11269] = 24'b010101010101010101010101;
rgb[11270] = 24'b011001100110011001100110;
rgb[11271] = 24'b011101110111011101110111;
rgb[11272] = 24'b100010001000100010001000;
rgb[11273] = 24'b100110011001100110011001;
rgb[11274] = 24'b101010101010101010101010;
rgb[11275] = 24'b101110111011101110111011;
rgb[11276] = 24'b110011001100110011001100;
rgb[11277] = 24'b110111011101110111011101;
rgb[11278] = 24'b111011101110111011101110;
rgb[11279] = 24'b111111111111111111111111;
rgb[11280] = 24'b000000000000000000000000;
rgb[11281] = 24'b000100000000111100010010;
rgb[11282] = 24'b001000000001111100100100;
rgb[11283] = 24'b001100000010111100110110;
rgb[11284] = 24'b010000010011111101001000;
rgb[11285] = 24'b010100010100111101011010;
rgb[11286] = 24'b011000010101111101101100;
rgb[11287] = 24'b011100100110111101111110;
rgb[11288] = 24'b100000111000000010001111;
rgb[11289] = 24'b100101001001001010011111;
rgb[11290] = 24'b101001101010010010101111;
rgb[11291] = 24'b101110001011011010111111;
rgb[11292] = 24'b110010011100100011001111;
rgb[11293] = 24'b110110111101101011011111;
rgb[11294] = 24'b111011011110110011101111;
rgb[11295] = 24'b111111111111111111111111;
rgb[11296] = 24'b000000000000000000000000;
rgb[11297] = 24'b000011110000111000010011;
rgb[11298] = 24'b000111110001110100100110;
rgb[11299] = 24'b001011100010110000111001;
rgb[11300] = 24'b001111100011101001001101;
rgb[11301] = 24'b010011010100100101100000;
rgb[11302] = 24'b010111010101100001110011;
rgb[11303] = 24'b011011010110011110000110;
rgb[11304] = 24'b011111100111100010010111;
rgb[11305] = 24'b100100001000101110100110;
rgb[11306] = 24'b101000101001111010110101;
rgb[11307] = 24'b101101011011000111000100;
rgb[11308] = 24'b110001111100010111010010;
rgb[11309] = 24'b110110101101100011100001;
rgb[11310] = 24'b111011001110101111110000;
rgb[11311] = 24'b111111111111111111111111;
rgb[11312] = 24'b000000000000000000000000;
rgb[11313] = 24'b000011100000110100010100;
rgb[11314] = 24'b000111010001101100101000;
rgb[11315] = 24'b001011000010100000111101;
rgb[11316] = 24'b001110110011011001010001;
rgb[11317] = 24'b010010100100010001100101;
rgb[11318] = 24'b010110010101000101111010;
rgb[11319] = 24'b011010000101111110001110;
rgb[11320] = 24'b011110010111000010011111;
rgb[11321] = 24'b100011001000010010101101;
rgb[11322] = 24'b100111111001100010111011;
rgb[11323] = 24'b101100101010110111001000;
rgb[11324] = 24'b110001011100000111010110;
rgb[11325] = 24'b110110001101011011100011;
rgb[11326] = 24'b111010111110101011110001;
rgb[11327] = 24'b111111111111111111111111;
rgb[11328] = 24'b000000000000000000000000;
rgb[11329] = 24'b000011100000110000010101;
rgb[11330] = 24'b000111000001100000101011;
rgb[11331] = 24'b001010100010010101000000;
rgb[11332] = 24'b001110000011000101010110;
rgb[11333] = 24'b010001100011111001101011;
rgb[11334] = 24'b010101010100101010000001;
rgb[11335] = 24'b011000110101011110010110;
rgb[11336] = 24'b011101000110100010100111;
rgb[11337] = 24'b100010000111110110110100;
rgb[11338] = 24'b100110111001001111000000;
rgb[11339] = 24'b101011111010100011001101;
rgb[11340] = 24'b110000111011111011011001;
rgb[11341] = 24'b110101111101001111100110;
rgb[11342] = 24'b111010111110100111110010;
rgb[11343] = 24'b111111111111111111111111;
rgb[11344] = 24'b000000000000000000000000;
rgb[11345] = 24'b000011010000101100010110;
rgb[11346] = 24'b000110100001011000101101;
rgb[11347] = 24'b001010000010001001000100;
rgb[11348] = 24'b001101010010110101011010;
rgb[11349] = 24'b010000110011100001110001;
rgb[11350] = 24'b010100000100010010001000;
rgb[11351] = 24'b010111100100111110011110;
rgb[11352] = 24'b011011110110000010101111;
rgb[11353] = 24'b100000110111011010111011;
rgb[11354] = 24'b100110001000110111000110;
rgb[11355] = 24'b101011001010010011010001;
rgb[11356] = 24'b110000011011101111011101;
rgb[11357] = 24'b110101011101000111101000;
rgb[11358] = 24'b111010101110100011110011;
rgb[11359] = 24'b111111111111111111111111;
rgb[11360] = 24'b000000000000000000000000;
rgb[11361] = 24'b000011000000101000010111;
rgb[11362] = 24'b000110010001010000101111;
rgb[11363] = 24'b001001100001111001000111;
rgb[11364] = 24'b001100110010100001011111;
rgb[11365] = 24'b001111110011001101110110;
rgb[11366] = 24'b010011000011110110001110;
rgb[11367] = 24'b010110010100011110100110;
rgb[11368] = 24'b011010100101100010110111;
rgb[11369] = 24'b011111110111000011000001;
rgb[11370] = 24'b100101001000011111001100;
rgb[11371] = 24'b101010101001111111010110;
rgb[11372] = 24'b101111111011011111100000;
rgb[11373] = 24'b110101001100111111101010;
rgb[11374] = 24'b111010011110011111110100;
rgb[11375] = 24'b111111111111111111111110;
rgb[11376] = 24'b000000000000000000000000;
rgb[11377] = 24'b000011000000100100011000;
rgb[11378] = 24'b000110000001001000110001;
rgb[11379] = 24'b001001000001101101001010;
rgb[11380] = 24'b001100000010010001100011;
rgb[11381] = 24'b001111000010110101111100;
rgb[11382] = 24'b010010000011011010010101;
rgb[11383] = 24'b010101000011111110101110;
rgb[11384] = 24'b011001010101000010111111;
rgb[11385] = 24'b011110110110100111001000;
rgb[11386] = 24'b100100011000001011010001;
rgb[11387] = 24'b101001111001101111011010;
rgb[11388] = 24'b101111011011010011100011;
rgb[11389] = 24'b110100111100110111101100;
rgb[11390] = 24'b111010011110011011110101;
rgb[11391] = 24'b111111111111111111111111;
rgb[11392] = 24'b000000000000000000000000;
rgb[11393] = 24'b000010110000011100011010;
rgb[11394] = 24'b000101100000111100110100;
rgb[11395] = 24'b001000100001011101001110;
rgb[11396] = 24'b001011010001111101101000;
rgb[11397] = 24'b001110000010011110000010;
rgb[11398] = 24'b010001000010111110011100;
rgb[11399] = 24'b010011110011011110110110;
rgb[11400] = 24'b011000000100100011000111;
rgb[11401] = 24'b011101110110001011001111;
rgb[11402] = 24'b100011010111110011010111;
rgb[11403] = 24'b101001001001011011011111;
rgb[11404] = 24'b101110111011000011100111;
rgb[11405] = 24'b110100011100101011101111;
rgb[11406] = 24'b111010001110010011110111;
rgb[11407] = 24'b111111111111111111111110;
rgb[11408] = 24'b000000000000000000000000;
rgb[11409] = 24'b000010100000011000011011;
rgb[11410] = 24'b000101010000110100110110;
rgb[11411] = 24'b001000000001010001010001;
rgb[11412] = 24'b001010100001101101101100;
rgb[11413] = 24'b001101010010000110001000;
rgb[11414] = 24'b010000000010100010100011;
rgb[11415] = 24'b010010100010111110111110;
rgb[11416] = 24'b010110110100000011001111;
rgb[11417] = 24'b011100110101101111010110;
rgb[11418] = 24'b100010100111011011011101;
rgb[11419] = 24'b101000011001001011100011;
rgb[11420] = 24'b101110011010110111101010;
rgb[11421] = 24'b110100001100100011110001;
rgb[11422] = 24'b111001111110001111111000;
rgb[11423] = 24'b111111111111111111111111;
rgb[11424] = 24'b000000000000000000000000;
rgb[11425] = 24'b000010010000010100011100;
rgb[11426] = 24'b000100110000101100111000;
rgb[11427] = 24'b000111010001000101010101;
rgb[11428] = 24'b001001110001011001110001;
rgb[11429] = 24'b001100010001110010001101;
rgb[11430] = 24'b001110110010001010101010;
rgb[11431] = 24'b010001010010011111000110;
rgb[11432] = 24'b010101100011100011010111;
rgb[11433] = 24'b011011100101010011011101;
rgb[11434] = 24'b100001100111000111100010;
rgb[11435] = 24'b100111101000110111101000;
rgb[11436] = 24'b101101101010101011101110;
rgb[11437] = 24'b110011101100011011110011;
rgb[11438] = 24'b111001101110001011111001;
rgb[11439] = 24'b111111111111111111111110;
rgb[11440] = 24'b000000000000000000000000;
rgb[11441] = 24'b000010010000010000011101;
rgb[11442] = 24'b000100100000100100111010;
rgb[11443] = 24'b000110110000110101011000;
rgb[11444] = 24'b001001010001001001110101;
rgb[11445] = 24'b001011100001011010010011;
rgb[11446] = 24'b001101110001101110110000;
rgb[11447] = 24'b010000000001111111001110;
rgb[11448] = 24'b010100010011000011011111;
rgb[11449] = 24'b011010100100111011100011;
rgb[11450] = 24'b100000110110101111101000;
rgb[11451] = 24'b100111001000100111101100;
rgb[11452] = 24'b101101001010011011110001;
rgb[11453] = 24'b110011011100010011110101;
rgb[11454] = 24'b111001101110000111111010;
rgb[11455] = 24'b111111111111111111111111;
rgb[11456] = 24'b000000000000000000000000;
rgb[11457] = 24'b000010000000001100011110;
rgb[11458] = 24'b000100010000011000111101;
rgb[11459] = 24'b000110010000101001011011;
rgb[11460] = 24'b001000100000110101111010;
rgb[11461] = 24'b001010100001000010011001;
rgb[11462] = 24'b001100110001010010110111;
rgb[11463] = 24'b001111000001011111010110;
rgb[11464] = 24'b010011010010100011100111;
rgb[11465] = 24'b011001100100011111101010;
rgb[11466] = 24'b011111110110010111101110;
rgb[11467] = 24'b100110011000010011110001;
rgb[11468] = 24'b101100101010001111110100;
rgb[11469] = 24'b110011001100000111111000;
rgb[11470] = 24'b111001011110000011111011;
rgb[11471] = 24'b111111111111111111111111;
rgb[11472] = 24'b000000000000000000000000;
rgb[11473] = 24'b000001110000001000011111;
rgb[11474] = 24'b000011110000010000111111;
rgb[11475] = 24'b000101110000011001011111;
rgb[11476] = 24'b000111110000100101111110;
rgb[11477] = 24'b001001110000101110011110;
rgb[11478] = 24'b001011110000110110111110;
rgb[11479] = 24'b001101110000111111011110;
rgb[11480] = 24'b010010000010000011101111;
rgb[11481] = 24'b011000100100000011110001;
rgb[11482] = 24'b011111000110000011110011;
rgb[11483] = 24'b100101101000000011110101;
rgb[11484] = 24'b101100001001111111111000;
rgb[11485] = 24'b110010101011111111111010;
rgb[11486] = 24'b111001001101111111111100;
rgb[11487] = 24'b111111111111111111111111;
rgb[11488] = 24'b000000000000000000000000;
rgb[11489] = 24'b000001110000000100100000;
rgb[11490] = 24'b000011100000001001000001;
rgb[11491] = 24'b000101010000001101100010;
rgb[11492] = 24'b000111000000010010000011;
rgb[11493] = 24'b001000110000010110100100;
rgb[11494] = 24'b001010110000011011000101;
rgb[11495] = 24'b001100100000011111100110;
rgb[11496] = 24'b010000110001100011110111;
rgb[11497] = 24'b010111100011100111111000;
rgb[11498] = 24'b011110000101101011111001;
rgb[11499] = 24'b100100110111101111111010;
rgb[11500] = 24'b101011101001110011111011;
rgb[11501] = 24'b110010011011110111111100;
rgb[11502] = 24'b111001001101111011111101;
rgb[11503] = 24'b111111111111111111111111;
rgb[11504] = 24'b000000000000000000000000;
rgb[11505] = 24'b000001100000000000100010;
rgb[11506] = 24'b000011000000000001000100;
rgb[11507] = 24'b000100110000000001100110;
rgb[11508] = 24'b000110010000000010001000;
rgb[11509] = 24'b001000000000000010101010;
rgb[11510] = 24'b001001100000000011001100;
rgb[11511] = 24'b001011010000000011101110;
rgb[11512] = 24'b001111100001000111111110;
rgb[11513] = 24'b010110010011001011111111;
rgb[11514] = 24'b011101010101010111111110;
rgb[11515] = 24'b100100000111011011111111;
rgb[11516] = 24'b101011001001100111111111;
rgb[11517] = 24'b110001111011101111111111;
rgb[11518] = 24'b111000111101110111111111;
rgb[11519] = 24'b111111111111111111111111;
rgb[11520] = 24'b000000000000000000000000;
rgb[11521] = 24'b000100010001000100010001;
rgb[11522] = 24'b001000100010001000100010;
rgb[11523] = 24'b001100110011001100110011;
rgb[11524] = 24'b010001000100010001000100;
rgb[11525] = 24'b010101010101010101010101;
rgb[11526] = 24'b011001100110011001100110;
rgb[11527] = 24'b011101110111011101110111;
rgb[11528] = 24'b100010001000100010001000;
rgb[11529] = 24'b100110011001100110011001;
rgb[11530] = 24'b101010101010101010101010;
rgb[11531] = 24'b101110111011101110111011;
rgb[11532] = 24'b110011001100110011001100;
rgb[11533] = 24'b110111011101110111011101;
rgb[11534] = 24'b111011101110111011101110;
rgb[11535] = 24'b111111111111111111111111;
rgb[11536] = 24'b000000000000000000000000;
rgb[11537] = 24'b000100000000111100010010;
rgb[11538] = 24'b001000010001111100100100;
rgb[11539] = 24'b001100010010111100110110;
rgb[11540] = 24'b010000100011111101001000;
rgb[11541] = 24'b010100100100111101011010;
rgb[11542] = 24'b011000110101111101101100;
rgb[11543] = 24'b011100110110111101111110;
rgb[11544] = 24'b100001001000000010001111;
rgb[11545] = 24'b100101101001001010011111;
rgb[11546] = 24'b101001111010010010101111;
rgb[11547] = 24'b101110011011011010111111;
rgb[11548] = 24'b110010101100100011001111;
rgb[11549] = 24'b110111001101101011011111;
rgb[11550] = 24'b111011011110110011101111;
rgb[11551] = 24'b111111111111111111111111;
rgb[11552] = 24'b000000000000000000000000;
rgb[11553] = 24'b000100000000111000010011;
rgb[11554] = 24'b001000000001110100100110;
rgb[11555] = 24'b001100000010110000111001;
rgb[11556] = 24'b010000000011101001001101;
rgb[11557] = 24'b010100000100100101100000;
rgb[11558] = 24'b011000000101100001110011;
rgb[11559] = 24'b011100000110011110000110;
rgb[11560] = 24'b100000010111100010010111;
rgb[11561] = 24'b100100111000101110100110;
rgb[11562] = 24'b101001011001111010110101;
rgb[11563] = 24'b101101111011000111000100;
rgb[11564] = 24'b110010011100010111010010;
rgb[11565] = 24'b110110111101100011100001;
rgb[11566] = 24'b111011011110101111110000;
rgb[11567] = 24'b111111111111111111111111;
rgb[11568] = 24'b000000000000000000000000;
rgb[11569] = 24'b000011110000110100010100;
rgb[11570] = 24'b000111110001101100101000;
rgb[11571] = 24'b001011100010100000111101;
rgb[11572] = 24'b001111100011011001010001;
rgb[11573] = 24'b010011010100010001100101;
rgb[11574] = 24'b010111010101000101111010;
rgb[11575] = 24'b011011000101111110001110;
rgb[11576] = 24'b011111010111000010011111;
rgb[11577] = 24'b100100001000010010101101;
rgb[11578] = 24'b101000101001100010111011;
rgb[11579] = 24'b101101011010110111001000;
rgb[11580] = 24'b110001111100000111010110;
rgb[11581] = 24'b110110101101011011100011;
rgb[11582] = 24'b111011001110101011110001;
rgb[11583] = 24'b111111111111111111111111;
rgb[11584] = 24'b000000000000000000000000;
rgb[11585] = 24'b000011110000110000010101;
rgb[11586] = 24'b000111100001100000101011;
rgb[11587] = 24'b001011010010010101000000;
rgb[11588] = 24'b001111000011000101010110;
rgb[11589] = 24'b010010110011111001101011;
rgb[11590] = 24'b010110100100101010000001;
rgb[11591] = 24'b011010010101011110010110;
rgb[11592] = 24'b011110100110100010100111;
rgb[11593] = 24'b100011010111110110110100;
rgb[11594] = 24'b101000001001001111000000;
rgb[11595] = 24'b101100111010100011001101;
rgb[11596] = 24'b110001101011111011011001;
rgb[11597] = 24'b110110011101001111100110;
rgb[11598] = 24'b111011001110100111110010;
rgb[11599] = 24'b111111111111111111111111;
rgb[11600] = 24'b000000000000000000000000;
rgb[11601] = 24'b000011100000101100010110;
rgb[11602] = 24'b000111010001011000101101;
rgb[11603] = 24'b001010110010001001000100;
rgb[11604] = 24'b001110100010110101011010;
rgb[11605] = 24'b010010000011100001110001;
rgb[11606] = 24'b010101110100010010001000;
rgb[11607] = 24'b011001100100111110011110;
rgb[11608] = 24'b011101110110000010101111;
rgb[11609] = 24'b100010100111011010111011;
rgb[11610] = 24'b100111011000110111000110;
rgb[11611] = 24'b101100011010010011010001;
rgb[11612] = 24'b110001001011101111011101;
rgb[11613] = 24'b110110001101000111101000;
rgb[11614] = 24'b111010111110100011110011;
rgb[11615] = 24'b111111111111111111111111;
rgb[11616] = 24'b000000000000000000000000;
rgb[11617] = 24'b000011100000101000010111;
rgb[11618] = 24'b000111000001010000101111;
rgb[11619] = 24'b001010100001111001000111;
rgb[11620] = 24'b001110000010100001011111;
rgb[11621] = 24'b010001100011001101110110;
rgb[11622] = 24'b010101000011110110001110;
rgb[11623] = 24'b011000100100011110100110;
rgb[11624] = 24'b011100110101100010110111;
rgb[11625] = 24'b100001110111000011000001;
rgb[11626] = 24'b100110111000011111001100;
rgb[11627] = 24'b101011111001111111010110;
rgb[11628] = 24'b110000111011011111100000;
rgb[11629] = 24'b110101111100111111101010;
rgb[11630] = 24'b111010111110011111110100;
rgb[11631] = 24'b111111111111111111111110;
rgb[11632] = 24'b000000000000000000000000;
rgb[11633] = 24'b000011010000100100011000;
rgb[11634] = 24'b000110110001001000110001;
rgb[11635] = 24'b001010000001101101001010;
rgb[11636] = 24'b001101100010010001100011;
rgb[11637] = 24'b010001000010110101111100;
rgb[11638] = 24'b010100010011011010010101;
rgb[11639] = 24'b010111110011111110101110;
rgb[11640] = 24'b011100000101000010111111;
rgb[11641] = 24'b100001000110100111001000;
rgb[11642] = 24'b100110011000001011010001;
rgb[11643] = 24'b101011011001101111011010;
rgb[11644] = 24'b110000011011010011100011;
rgb[11645] = 24'b110101101100110111101100;
rgb[11646] = 24'b111010101110011011110101;
rgb[11647] = 24'b111111111111111111111111;
rgb[11648] = 24'b000000000000000000000000;
rgb[11649] = 24'b000011010000011100011010;
rgb[11650] = 24'b000110100000111100110100;
rgb[11651] = 24'b001001110001011101001110;
rgb[11652] = 24'b001101000001111101101000;
rgb[11653] = 24'b010000010010011110000010;
rgb[11654] = 24'b010011100010111110011100;
rgb[11655] = 24'b010110110011011110110110;
rgb[11656] = 24'b011011000100100011000111;
rgb[11657] = 24'b100000010110001011001111;
rgb[11658] = 24'b100101100111110011010111;
rgb[11659] = 24'b101010111001011011011111;
rgb[11660] = 24'b110000001011000011100111;
rgb[11661] = 24'b110101011100101011101111;
rgb[11662] = 24'b111010101110010011110111;
rgb[11663] = 24'b111111111111111111111110;
rgb[11664] = 24'b000000000000000000000000;
rgb[11665] = 24'b000011000000011000011011;
rgb[11666] = 24'b000110010000110100110110;
rgb[11667] = 24'b001001010001010001010001;
rgb[11668] = 24'b001100100001101101101100;
rgb[11669] = 24'b001111110010000110001000;
rgb[11670] = 24'b010010110010100010100011;
rgb[11671] = 24'b010110000010111110111110;
rgb[11672] = 24'b011010010100000011001111;
rgb[11673] = 24'b011111100101101111010110;
rgb[11674] = 24'b100101000111011011011101;
rgb[11675] = 24'b101010011001001011100011;
rgb[11676] = 24'b101111101010110111101010;
rgb[11677] = 24'b110101001100100011110001;
rgb[11678] = 24'b111010011110001111111000;
rgb[11679] = 24'b111111111111111111111111;
rgb[11680] = 24'b000000000000000000000000;
rgb[11681] = 24'b000011000000010100011100;
rgb[11682] = 24'b000110000000101100111000;
rgb[11683] = 24'b001001000001000101010101;
rgb[11684] = 24'b001100000001011001110001;
rgb[11685] = 24'b001111000001110010001101;
rgb[11686] = 24'b010010000010001010101010;
rgb[11687] = 24'b010101010010011111000110;
rgb[11688] = 24'b011001100011100011010111;
rgb[11689] = 24'b011110110101010011011101;
rgb[11690] = 24'b100100010111000111100010;
rgb[11691] = 24'b101001111000110111101000;
rgb[11692] = 24'b101111011010101011101110;
rgb[11693] = 24'b110100111100011011110011;
rgb[11694] = 24'b111010011110001011111001;
rgb[11695] = 24'b111111111111111111111110;
rgb[11696] = 24'b000000000000000000000000;
rgb[11697] = 24'b000010110000010000011101;
rgb[11698] = 24'b000101110000100100111010;
rgb[11699] = 24'b001000100000110101011000;
rgb[11700] = 24'b001011100001001001110101;
rgb[11701] = 24'b001110100001011010010011;
rgb[11702] = 24'b010001010001101110110000;
rgb[11703] = 24'b010100010001111111001110;
rgb[11704] = 24'b011000100011000011011111;
rgb[11705] = 24'b011110000100111011100011;
rgb[11706] = 24'b100011110110101111101000;
rgb[11707] = 24'b101001011000100111101100;
rgb[11708] = 24'b101110111010011011110001;
rgb[11709] = 24'b110100101100010011110101;
rgb[11710] = 24'b111010001110000111111010;
rgb[11711] = 24'b111111111111111111111111;
rgb[11712] = 24'b000000000000000000000000;
rgb[11713] = 24'b000010110000001100011110;
rgb[11714] = 24'b000101100000011000111101;
rgb[11715] = 24'b001000010000101001011011;
rgb[11716] = 24'b001011000000110101111010;
rgb[11717] = 24'b001101110001000010011001;
rgb[11718] = 24'b010000110001010010110111;
rgb[11719] = 24'b010011100001011111010110;
rgb[11720] = 24'b010111110010100011100111;
rgb[11721] = 24'b011101100100011111101010;
rgb[11722] = 24'b100011000110010111101110;
rgb[11723] = 24'b101000111000010011110001;
rgb[11724] = 24'b101110101010001111110100;
rgb[11725] = 24'b110100011100000111111000;
rgb[11726] = 24'b111010001110000011111011;
rgb[11727] = 24'b111111111111111111111111;
rgb[11728] = 24'b000000000000000000000000;
rgb[11729] = 24'b000010100000001000011111;
rgb[11730] = 24'b000101010000010000111111;
rgb[11731] = 24'b001000000000011001011111;
rgb[11732] = 24'b001010100000100101111110;
rgb[11733] = 24'b001101010000101110011110;
rgb[11734] = 24'b010000000000110110111110;
rgb[11735] = 24'b010010100000111111011110;
rgb[11736] = 24'b010110110010000011101111;
rgb[11737] = 24'b011100110100000011110001;
rgb[11738] = 24'b100010100110000011110011;
rgb[11739] = 24'b101000011000000011110101;
rgb[11740] = 24'b101110011001111111111000;
rgb[11741] = 24'b110100001011111111111010;
rgb[11742] = 24'b111001111101111111111100;
rgb[11743] = 24'b111111111111111111111111;
rgb[11744] = 24'b000000000000000000000000;
rgb[11745] = 24'b000010100000000100100000;
rgb[11746] = 24'b000101000000001001000001;
rgb[11747] = 24'b000111100000001101100010;
rgb[11748] = 24'b001010000000010010000011;
rgb[11749] = 24'b001100110000010110100100;
rgb[11750] = 24'b001111010000011011000101;
rgb[11751] = 24'b010001110000011111100110;
rgb[11752] = 24'b010110000001100011110111;
rgb[11753] = 24'b011100000011100111111000;
rgb[11754] = 24'b100010000101101011111001;
rgb[11755] = 24'b100111110111101111111010;
rgb[11756] = 24'b101101111001110011111011;
rgb[11757] = 24'b110011111011110111111100;
rgb[11758] = 24'b111001111101111011111101;
rgb[11759] = 24'b111111111111111111111111;
rgb[11760] = 24'b000000000000000000000000;
rgb[11761] = 24'b000010010000000000100010;
rgb[11762] = 24'b000100110000000001000100;
rgb[11763] = 24'b000111010000000001100110;
rgb[11764] = 24'b001001100000000010001000;
rgb[11765] = 24'b001100000000000010101010;
rgb[11766] = 24'b001110100000000011001100;
rgb[11767] = 24'b010001000000000011101110;
rgb[11768] = 24'b010101010001000111111110;
rgb[11769] = 24'b011011010011001011111111;
rgb[11770] = 24'b100001010101010111111110;
rgb[11771] = 24'b100111010111011011111111;
rgb[11772] = 24'b101101101001100111111111;
rgb[11773] = 24'b110011101011101111111111;
rgb[11774] = 24'b111001101101110111111111;
rgb[11775] = 24'b111111111111111111111111;
rgb[11776] = 24'b000000000000000000000000;
rgb[11777] = 24'b000100010001000100010001;
rgb[11778] = 24'b001000100010001000100010;
rgb[11779] = 24'b001100110011001100110011;
rgb[11780] = 24'b010001000100010001000100;
rgb[11781] = 24'b010101010101010101010101;
rgb[11782] = 24'b011001100110011001100110;
rgb[11783] = 24'b011101110111011101110111;
rgb[11784] = 24'b100010001000100010001000;
rgb[11785] = 24'b100110011001100110011001;
rgb[11786] = 24'b101010101010101010101010;
rgb[11787] = 24'b101110111011101110111011;
rgb[11788] = 24'b110011001100110011001100;
rgb[11789] = 24'b110111011101110111011101;
rgb[11790] = 24'b111011101110111011101110;
rgb[11791] = 24'b111111111111111111111111;
rgb[11792] = 24'b000000000000000000000000;
rgb[11793] = 24'b000100000000111100010010;
rgb[11794] = 24'b001000010001111100100100;
rgb[11795] = 24'b001100100010111100110110;
rgb[11796] = 24'b010000100011111101001000;
rgb[11797] = 24'b010100110100111101011010;
rgb[11798] = 24'b011001000101111101101100;
rgb[11799] = 24'b011101010110111101111110;
rgb[11800] = 24'b100001101000000010001111;
rgb[11801] = 24'b100101111001001010011111;
rgb[11802] = 24'b101010001010010010101111;
rgb[11803] = 24'b101110011011011010111111;
rgb[11804] = 24'b110010111100100011001111;
rgb[11805] = 24'b110111001101101011011111;
rgb[11806] = 24'b111011011110110011101111;
rgb[11807] = 24'b111111111111111111111111;
rgb[11808] = 24'b000000000000000000000000;
rgb[11809] = 24'b000100000000111000010011;
rgb[11810] = 24'b001000000001110100100110;
rgb[11811] = 24'b001100010010110000111001;
rgb[11812] = 24'b010000010011101001001101;
rgb[11813] = 24'b010100100100100101100000;
rgb[11814] = 24'b011000100101100001110011;
rgb[11815] = 24'b011100110110011110000110;
rgb[11816] = 24'b100001000111100010010111;
rgb[11817] = 24'b100101011000101110100110;
rgb[11818] = 24'b101001111001111010110101;
rgb[11819] = 24'b101110001011000111000100;
rgb[11820] = 24'b110010101100010111010010;
rgb[11821] = 24'b110110111101100011100001;
rgb[11822] = 24'b111011011110101111110000;
rgb[11823] = 24'b111111111111111111111111;
rgb[11824] = 24'b000000000000000000000000;
rgb[11825] = 24'b000100000000110100010100;
rgb[11826] = 24'b001000000001101100101000;
rgb[11827] = 24'b001100000010100000111101;
rgb[11828] = 24'b010000000011011001010001;
rgb[11829] = 24'b010100000100010001100101;
rgb[11830] = 24'b011000010101000101111010;
rgb[11831] = 24'b011100010101111110001110;
rgb[11832] = 24'b100000100111000010011111;
rgb[11833] = 24'b100101001000010010101101;
rgb[11834] = 24'b101001011001100010111011;
rgb[11835] = 24'b101101111010110111001000;
rgb[11836] = 24'b110010011100000111010110;
rgb[11837] = 24'b110110111101011011100011;
rgb[11838] = 24'b111011011110101011110001;
rgb[11839] = 24'b111111111111111111111111;
rgb[11840] = 24'b000000000000000000000000;
rgb[11841] = 24'b000011110000110000010101;
rgb[11842] = 24'b000111110001100000101011;
rgb[11843] = 24'b001011110010010101000000;
rgb[11844] = 24'b001111110011000101010110;
rgb[11845] = 24'b010011110011111001101011;
rgb[11846] = 24'b010111110100101010000001;
rgb[11847] = 24'b011011110101011110010110;
rgb[11848] = 24'b100000000110100010100111;
rgb[11849] = 24'b100100100111110110110100;
rgb[11850] = 24'b101001001001001111000000;
rgb[11851] = 24'b101101101010100011001101;
rgb[11852] = 24'b110010001011111011011001;
rgb[11853] = 24'b110110101101001111100110;
rgb[11854] = 24'b111011001110100111110010;
rgb[11855] = 24'b111111111111111111111111;
rgb[11856] = 24'b000000000000000000000000;
rgb[11857] = 24'b000011110000101100010110;
rgb[11858] = 24'b000111110001011000101101;
rgb[11859] = 24'b001011100010001001000100;
rgb[11860] = 24'b001111100010110101011010;
rgb[11861] = 24'b010011100011100001110001;
rgb[11862] = 24'b010111010100010010001000;
rgb[11863] = 24'b011011010100111110011110;
rgb[11864] = 24'b011111100110000010101111;
rgb[11865] = 24'b100100000111011010111011;
rgb[11866] = 24'b101000111000110111000110;
rgb[11867] = 24'b101101011010010011010001;
rgb[11868] = 24'b110001111011101111011101;
rgb[11869] = 24'b110110101101000111101000;
rgb[11870] = 24'b111011001110100011110011;
rgb[11871] = 24'b111111111111111111111111;
rgb[11872] = 24'b000000000000000000000000;
rgb[11873] = 24'b000011110000101000010111;
rgb[11874] = 24'b000111100001010000101111;
rgb[11875] = 24'b001011100001111001000111;
rgb[11876] = 24'b001111010010100001011111;
rgb[11877] = 24'b010011000011001101110110;
rgb[11878] = 24'b010111000011110110001110;
rgb[11879] = 24'b011010110100011110100110;
rgb[11880] = 24'b011111000101100010110111;
rgb[11881] = 24'b100011110111000011000001;
rgb[11882] = 24'b101000011000011111001100;
rgb[11883] = 24'b101101001001111111010110;
rgb[11884] = 24'b110001111011011111100000;
rgb[11885] = 24'b110110011100111111101010;
rgb[11886] = 24'b111011001110011111110100;
rgb[11887] = 24'b111111111111111111111110;
rgb[11888] = 24'b000000000000000000000000;
rgb[11889] = 24'b000011110000100100011000;
rgb[11890] = 24'b000111100001001000110001;
rgb[11891] = 24'b001011010001101101001010;
rgb[11892] = 24'b001111000010010001100011;
rgb[11893] = 24'b010010110010110101111100;
rgb[11894] = 24'b010110100011011010010101;
rgb[11895] = 24'b011010010011111110101110;
rgb[11896] = 24'b011110100101000010111111;
rgb[11897] = 24'b100011010110100111001000;
rgb[11898] = 24'b101000001000001011010001;
rgb[11899] = 24'b101100111001101111011010;
rgb[11900] = 24'b110001101011010011100011;
rgb[11901] = 24'b110110011100110111101100;
rgb[11902] = 24'b111011001110011011110101;
rgb[11903] = 24'b111111111111111111111111;
rgb[11904] = 24'b000000000000000000000000;
rgb[11905] = 24'b000011100000011100011010;
rgb[11906] = 24'b000111010000111100110100;
rgb[11907] = 24'b001011000001011101001110;
rgb[11908] = 24'b001110110001111101101000;
rgb[11909] = 24'b010010100010011110000010;
rgb[11910] = 24'b010110010010111110011100;
rgb[11911] = 24'b011001110011011110110110;
rgb[11912] = 24'b011110000100100011000111;
rgb[11913] = 24'b100011000110001011001111;
rgb[11914] = 24'b100111110111110011010111;
rgb[11915] = 24'b101100101001011011011111;
rgb[11916] = 24'b110001011011000011100111;
rgb[11917] = 24'b110110001100101011101111;
rgb[11918] = 24'b111010111110010011110111;
rgb[11919] = 24'b111111111111111111111110;
rgb[11920] = 24'b000000000000000000000000;
rgb[11921] = 24'b000011100000011000011011;
rgb[11922] = 24'b000111010000110100110110;
rgb[11923] = 24'b001010110001010001010001;
rgb[11924] = 24'b001110100001101101101100;
rgb[11925] = 24'b010010000010000110001000;
rgb[11926] = 24'b010101110010100010100011;
rgb[11927] = 24'b011001010010111110111110;
rgb[11928] = 24'b011101110100000011001111;
rgb[11929] = 24'b100010100101101111010110;
rgb[11930] = 24'b100111010111011011011101;
rgb[11931] = 24'b101100011001001011100011;
rgb[11932] = 24'b110001001010110111101010;
rgb[11933] = 24'b110110001100100011110001;
rgb[11934] = 24'b111010111110001111111000;
rgb[11935] = 24'b111111111111111111111111;
rgb[11936] = 24'b000000000000000000000000;
rgb[11937] = 24'b000011100000010100011100;
rgb[11938] = 24'b000111000000101100111000;
rgb[11939] = 24'b001010100001000101010101;
rgb[11940] = 24'b001110010001011001110001;
rgb[11941] = 24'b010001110001110010001101;
rgb[11942] = 24'b010101010010001010101010;
rgb[11943] = 24'b011001000010011111000110;
rgb[11944] = 24'b011101010011100011010111;
rgb[11945] = 24'b100010000101010011011101;
rgb[11946] = 24'b100111000111000111100010;
rgb[11947] = 24'b101100001000110111101000;
rgb[11948] = 24'b110000111010101011101110;
rgb[11949] = 24'b110101111100011011110011;
rgb[11950] = 24'b111010111110001011111001;
rgb[11951] = 24'b111111111111111111111110;
rgb[11952] = 24'b000000000000000000000000;
rgb[11953] = 24'b000011100000010000011101;
rgb[11954] = 24'b000111000000100100111010;
rgb[11955] = 24'b001010100000110101011000;
rgb[11956] = 24'b001110000001001001110101;
rgb[11957] = 24'b010001100001011010010011;
rgb[11958] = 24'b010101000001101110110000;
rgb[11959] = 24'b011000100001111111001110;
rgb[11960] = 24'b011100110011000011011111;
rgb[11961] = 24'b100001110100111011100011;
rgb[11962] = 24'b100110110110101111101000;
rgb[11963] = 24'b101011111000100111101100;
rgb[11964] = 24'b110000111010011011110001;
rgb[11965] = 24'b110101111100010011110101;
rgb[11966] = 24'b111010111110000111111010;
rgb[11967] = 24'b111111111111111111111111;
rgb[11968] = 24'b000000000000000000000000;
rgb[11969] = 24'b000011010000001100011110;
rgb[11970] = 24'b000110110000011000111101;
rgb[11971] = 24'b001010010000101001011011;
rgb[11972] = 24'b001101110000110101111010;
rgb[11973] = 24'b010001000001000010011001;
rgb[11974] = 24'b010100100001010010110111;
rgb[11975] = 24'b011000000001011111010110;
rgb[11976] = 24'b011100010010100011100111;
rgb[11977] = 24'b100001010100011111101010;
rgb[11978] = 24'b100110010110010111101110;
rgb[11979] = 24'b101011101000010011110001;
rgb[11980] = 24'b110000101010001111110100;
rgb[11981] = 24'b110101101100000111111000;
rgb[11982] = 24'b111010101110000011111011;
rgb[11983] = 24'b111111111111111111111111;
rgb[11984] = 24'b000000000000000000000000;
rgb[11985] = 24'b000011010000001000011111;
rgb[11986] = 24'b000110100000010000111111;
rgb[11987] = 24'b001010000000011001011111;
rgb[11988] = 24'b001101010000100101111110;
rgb[11989] = 24'b010000110000101110011110;
rgb[11990] = 24'b010100000000110110111110;
rgb[11991] = 24'b010111100000111111011110;
rgb[11992] = 24'b011011110010000011101111;
rgb[11993] = 24'b100000110100000011110001;
rgb[11994] = 24'b100110000110000011110011;
rgb[11995] = 24'b101011001000000011110101;
rgb[11996] = 24'b110000011001111111111000;
rgb[11997] = 24'b110101011011111111111010;
rgb[11998] = 24'b111010101101111111111100;
rgb[11999] = 24'b111111111111111111111111;
rgb[12000] = 24'b000000000000000000000000;
rgb[12001] = 24'b000011010000000100100000;
rgb[12002] = 24'b000110100000001001000001;
rgb[12003] = 24'b001001110000001101100010;
rgb[12004] = 24'b001101000000010010000011;
rgb[12005] = 24'b010000100000010110100100;
rgb[12006] = 24'b010011110000011011000101;
rgb[12007] = 24'b010111000000011111100110;
rgb[12008] = 24'b011011010001100011110111;
rgb[12009] = 24'b100000100011100111111000;
rgb[12010] = 24'b100101110101101011111001;
rgb[12011] = 24'b101010110111101111111010;
rgb[12012] = 24'b110000001001110011111011;
rgb[12013] = 24'b110101011011110111111100;
rgb[12014] = 24'b111010101101111011111101;
rgb[12015] = 24'b111111111111111111111111;
rgb[12016] = 24'b000000000000000000000000;
rgb[12017] = 24'b000011000000000000100010;
rgb[12018] = 24'b000110010000000001000100;
rgb[12019] = 24'b001001100000000001100110;
rgb[12020] = 24'b001100110000000010001000;
rgb[12021] = 24'b010000000000000010101010;
rgb[12022] = 24'b010011010000000011001100;
rgb[12023] = 24'b010110100000000011101110;
rgb[12024] = 24'b011010110001000111111110;
rgb[12025] = 24'b100000000011001011111111;
rgb[12026] = 24'b100101010101010111111110;
rgb[12027] = 24'b101010100111011011111111;
rgb[12028] = 24'b101111111001100111111111;
rgb[12029] = 24'b110101001011101111111111;
rgb[12030] = 24'b111010011101110111111111;
rgb[12031] = 24'b111111111111111111111111;
rgb[12032] = 24'b000000000000000000000000;
rgb[12033] = 24'b000100010001000100010001;
rgb[12034] = 24'b001000100010001000100010;
rgb[12035] = 24'b001100110011001100110011;
rgb[12036] = 24'b010001000100010001000100;
rgb[12037] = 24'b010101010101010101010101;
rgb[12038] = 24'b011001100110011001100110;
rgb[12039] = 24'b011101110111011101110111;
rgb[12040] = 24'b100010001000100010001000;
rgb[12041] = 24'b100110011001100110011001;
rgb[12042] = 24'b101010101010101010101010;
rgb[12043] = 24'b101110111011101110111011;
rgb[12044] = 24'b110011001100110011001100;
rgb[12045] = 24'b110111011101110111011101;
rgb[12046] = 24'b111011101110111011101110;
rgb[12047] = 24'b111111111111111111111111;
rgb[12048] = 24'b000000000000000000000000;
rgb[12049] = 24'b000100000000111100010010;
rgb[12050] = 24'b001000010001111100100100;
rgb[12051] = 24'b001100100010111100110110;
rgb[12052] = 24'b010000110011111101001000;
rgb[12053] = 24'b010101000100111101011010;
rgb[12054] = 24'b011001010101111101101100;
rgb[12055] = 24'b011101100110111101111110;
rgb[12056] = 24'b100001111000000010001111;
rgb[12057] = 24'b100110001001001010011111;
rgb[12058] = 24'b101010011010010010101111;
rgb[12059] = 24'b101110101011011010111111;
rgb[12060] = 24'b110010111100100011001111;
rgb[12061] = 24'b110111001101101011011111;
rgb[12062] = 24'b111011011110110011101111;
rgb[12063] = 24'b111111111111111111111111;
rgb[12064] = 24'b000000000000000000000000;
rgb[12065] = 24'b000100000000111000010011;
rgb[12066] = 24'b001000010001110100100110;
rgb[12067] = 24'b001100100010110000111001;
rgb[12068] = 24'b010000110011101001001101;
rgb[12069] = 24'b010101000100100101100000;
rgb[12070] = 24'b011001010101100001110011;
rgb[12071] = 24'b011101100110011110000110;
rgb[12072] = 24'b100001110111100010010111;
rgb[12073] = 24'b100110001000101110100110;
rgb[12074] = 24'b101010011001111010110101;
rgb[12075] = 24'b101110101011000111000100;
rgb[12076] = 24'b110010111100010111010010;
rgb[12077] = 24'b110111001101100011100001;
rgb[12078] = 24'b111011011110101111110000;
rgb[12079] = 24'b111111111111111111111111;
rgb[12080] = 24'b000000000000000000000000;
rgb[12081] = 24'b000100000000110100010100;
rgb[12082] = 24'b001000010001101100101000;
rgb[12083] = 24'b001100100010100000111101;
rgb[12084] = 24'b010000110011011001010001;
rgb[12085] = 24'b010101000100010001100101;
rgb[12086] = 24'b011001010101000101111010;
rgb[12087] = 24'b011101010101111110001110;
rgb[12088] = 24'b100001100111000010011111;
rgb[12089] = 24'b100110001000010010101101;
rgb[12090] = 24'b101010011001100010111011;
rgb[12091] = 24'b101110101010110111001000;
rgb[12092] = 24'b110010111100000111010110;
rgb[12093] = 24'b110111001101011011100011;
rgb[12094] = 24'b111011011110101011110001;
rgb[12095] = 24'b111111111111111111111111;
rgb[12096] = 24'b000000000000000000000000;
rgb[12097] = 24'b000100000000110000010101;
rgb[12098] = 24'b001000010001100000101011;
rgb[12099] = 24'b001100100010010101000000;
rgb[12100] = 24'b010000110011000101010110;
rgb[12101] = 24'b010100110011111001101011;
rgb[12102] = 24'b011001000100101010000001;
rgb[12103] = 24'b011101010101011110010110;
rgb[12104] = 24'b100001100110100010100111;
rgb[12105] = 24'b100101110111110110110100;
rgb[12106] = 24'b101010001001001111000000;
rgb[12107] = 24'b101110101010100011001101;
rgb[12108] = 24'b110010111011111011011001;
rgb[12109] = 24'b110111001101001111100110;
rgb[12110] = 24'b111011011110100111110010;
rgb[12111] = 24'b111111111111111111111111;
rgb[12112] = 24'b000000000000000000000000;
rgb[12113] = 24'b000100000000101100010110;
rgb[12114] = 24'b001000010001011000101101;
rgb[12115] = 24'b001100100010001001000100;
rgb[12116] = 24'b010000100010110101011010;
rgb[12117] = 24'b010100110011100001110001;
rgb[12118] = 24'b011001000100010010001000;
rgb[12119] = 24'b011101010100111110011110;
rgb[12120] = 24'b100001100110000010101111;
rgb[12121] = 24'b100101110111011010111011;
rgb[12122] = 24'b101010001000110111000110;
rgb[12123] = 24'b101110011010010011010001;
rgb[12124] = 24'b110010111011101111011101;
rgb[12125] = 24'b110111001101000111101000;
rgb[12126] = 24'b111011011110100011110011;
rgb[12127] = 24'b111111111111111111111111;
rgb[12128] = 24'b000000000000000000000000;
rgb[12129] = 24'b000100000000101000010111;
rgb[12130] = 24'b001000010001010000101111;
rgb[12131] = 24'b001100100001111001000111;
rgb[12132] = 24'b010000100010100001011111;
rgb[12133] = 24'b010100110011001101110110;
rgb[12134] = 24'b011001000011110110001110;
rgb[12135] = 24'b011101000100011110100110;
rgb[12136] = 24'b100001010101100010110111;
rgb[12137] = 24'b100101110111000011000001;
rgb[12138] = 24'b101010001000011111001100;
rgb[12139] = 24'b101110011001111111010110;
rgb[12140] = 24'b110010111011011111100000;
rgb[12141] = 24'b110111001100111111101010;
rgb[12142] = 24'b111011011110011111110100;
rgb[12143] = 24'b111111111111111111111110;
rgb[12144] = 24'b000000000000000000000000;
rgb[12145] = 24'b000100000000100100011000;
rgb[12146] = 24'b001000010001001000110001;
rgb[12147] = 24'b001100010001101101001010;
rgb[12148] = 24'b010000100010010001100011;
rgb[12149] = 24'b010100110010110101111100;
rgb[12150] = 24'b011000110011011010010101;
rgb[12151] = 24'b011101000011111110101110;
rgb[12152] = 24'b100001010101000010111111;
rgb[12153] = 24'b100101100110100111001000;
rgb[12154] = 24'b101010001000001011010001;
rgb[12155] = 24'b101110011001101111011010;
rgb[12156] = 24'b110010101011010011100011;
rgb[12157] = 24'b110111001100110111101100;
rgb[12158] = 24'b111011011110011011110101;
rgb[12159] = 24'b111111111111111111111111;
rgb[12160] = 24'b000000000000000000000000;
rgb[12161] = 24'b000100000000011100011010;
rgb[12162] = 24'b001000010000111100110100;
rgb[12163] = 24'b001100010001011101001110;
rgb[12164] = 24'b010000100001111101101000;
rgb[12165] = 24'b010100100010011110000010;
rgb[12166] = 24'b011000110010111110011100;
rgb[12167] = 24'b011100110011011110110110;
rgb[12168] = 24'b100001000100100011000111;
rgb[12169] = 24'b100101100110001011001111;
rgb[12170] = 24'b101001110111110011010111;
rgb[12171] = 24'b101110011001011011011111;
rgb[12172] = 24'b110010101011000011100111;
rgb[12173] = 24'b110111001100101011101111;
rgb[12174] = 24'b111011011110010011110111;
rgb[12175] = 24'b111111111111111111111110;
rgb[12176] = 24'b000000000000000000000000;
rgb[12177] = 24'b000100000000011000011011;
rgb[12178] = 24'b001000010000110100110110;
rgb[12179] = 24'b001100010001010001010001;
rgb[12180] = 24'b010000100001101101101100;
rgb[12181] = 24'b010100100010000110001000;
rgb[12182] = 24'b011000110010100010100011;
rgb[12183] = 24'b011100110010111110111110;
rgb[12184] = 24'b100001000100000011001111;
rgb[12185] = 24'b100101100101101111010110;
rgb[12186] = 24'b101001110111011011011101;
rgb[12187] = 24'b101110011001001011100011;
rgb[12188] = 24'b110010101010110111101010;
rgb[12189] = 24'b110111001100100011110001;
rgb[12190] = 24'b111011011110001111111000;
rgb[12191] = 24'b111111111111111111111111;
rgb[12192] = 24'b000000000000000000000000;
rgb[12193] = 24'b000100000000010100011100;
rgb[12194] = 24'b001000000000101100111000;
rgb[12195] = 24'b001100010001000101010101;
rgb[12196] = 24'b010000010001011001110001;
rgb[12197] = 24'b010100100001110010001101;
rgb[12198] = 24'b011000100010001010101010;
rgb[12199] = 24'b011100110010011111000110;
rgb[12200] = 24'b100001000011100011010111;
rgb[12201] = 24'b100101010101010011011101;
rgb[12202] = 24'b101001110111000111100010;
rgb[12203] = 24'b101110001000110111101000;
rgb[12204] = 24'b110010101010101011101110;
rgb[12205] = 24'b110110111100011011110011;
rgb[12206] = 24'b111011011110001011111001;
rgb[12207] = 24'b111111111111111111111110;
rgb[12208] = 24'b000000000000000000000000;
rgb[12209] = 24'b000100000000010000011101;
rgb[12210] = 24'b001000000000100100111010;
rgb[12211] = 24'b001100010000110101011000;
rgb[12212] = 24'b010000010001001001110101;
rgb[12213] = 24'b010100100001011010010011;
rgb[12214] = 24'b011000100001101110110000;
rgb[12215] = 24'b011100100001111111001110;
rgb[12216] = 24'b100000110011000011011111;
rgb[12217] = 24'b100101010100111011100011;
rgb[12218] = 24'b101001110110101111101000;
rgb[12219] = 24'b101110001000100111101100;
rgb[12220] = 24'b110010101010011011110001;
rgb[12221] = 24'b110110111100010011110101;
rgb[12222] = 24'b111011011110000111111010;
rgb[12223] = 24'b111111111111111111111111;
rgb[12224] = 24'b000000000000000000000000;
rgb[12225] = 24'b000100000000001100011110;
rgb[12226] = 24'b001000000000011000111101;
rgb[12227] = 24'b001100010000101001011011;
rgb[12228] = 24'b010000010000110101111010;
rgb[12229] = 24'b010100010001000010011001;
rgb[12230] = 24'b011000100001010010110111;
rgb[12231] = 24'b011100100001011111010110;
rgb[12232] = 24'b100000110010100011100111;
rgb[12233] = 24'b100101010100011111101010;
rgb[12234] = 24'b101001100110010111101110;
rgb[12235] = 24'b101110001000010011110001;
rgb[12236] = 24'b110010101010001111110100;
rgb[12237] = 24'b110110111100000111111000;
rgb[12238] = 24'b111011011110000011111011;
rgb[12239] = 24'b111111111111111111111111;
rgb[12240] = 24'b000000000000000000000000;
rgb[12241] = 24'b000100000000001000011111;
rgb[12242] = 24'b001000000000010000111111;
rgb[12243] = 24'b001100000000011001011111;
rgb[12244] = 24'b010000010000100101111110;
rgb[12245] = 24'b010100010000101110011110;
rgb[12246] = 24'b011000010000110110111110;
rgb[12247] = 24'b011100100000111111011110;
rgb[12248] = 24'b100000110010000011101111;
rgb[12249] = 24'b100101000100000011110001;
rgb[12250] = 24'b101001100110000011110011;
rgb[12251] = 24'b101110001000000011110101;
rgb[12252] = 24'b110010011001111111111000;
rgb[12253] = 24'b110110111011111111111010;
rgb[12254] = 24'b111011011101111111111100;
rgb[12255] = 24'b111111111111111111111111;
rgb[12256] = 24'b000000000000000000000000;
rgb[12257] = 24'b000100000000000100100000;
rgb[12258] = 24'b001000000000001001000001;
rgb[12259] = 24'b001100000000001101100010;
rgb[12260] = 24'b010000000000010010000011;
rgb[12261] = 24'b010100010000010110100100;
rgb[12262] = 24'b011000010000011011000101;
rgb[12263] = 24'b011100010000011111100110;
rgb[12264] = 24'b100000100001100011110111;
rgb[12265] = 24'b100101000011100111111000;
rgb[12266] = 24'b101001100101101011111001;
rgb[12267] = 24'b101101110111101111111010;
rgb[12268] = 24'b110010011001110011111011;
rgb[12269] = 24'b110110111011110111111100;
rgb[12270] = 24'b111011011101111011111101;
rgb[12271] = 24'b111111111111111111111111;
rgb[12272] = 24'b000000000000000000000000;
rgb[12273] = 24'b000100000000000000100010;
rgb[12274] = 24'b001000000000000001000100;
rgb[12275] = 24'b001100000000000001100110;
rgb[12276] = 24'b010000000000000010001000;
rgb[12277] = 24'b010100000000000010101010;
rgb[12278] = 24'b011000010000000011001100;
rgb[12279] = 24'b011100010000000011101110;
rgb[12280] = 24'b100000100001000111111110;
rgb[12281] = 24'b100101000011001011111111;
rgb[12282] = 24'b101001010101010111111110;
rgb[12283] = 24'b101101110111011011111111;
rgb[12284] = 24'b110010011001100111111111;
rgb[12285] = 24'b110110111011101111111111;
rgb[12286] = 24'b111011011101110111111111;
rgb[12287] = 24'b111111111111111111111111;
rgb[12288] = 24'b000000000000000000000000;
rgb[12289] = 24'b000100010001000100010001;
rgb[12290] = 24'b001000100010001000100010;
rgb[12291] = 24'b001100110011001100110011;
rgb[12292] = 24'b010001000100010001000100;
rgb[12293] = 24'b010101010101010101010101;
rgb[12294] = 24'b011001100110011001100110;
rgb[12295] = 24'b011101110111011101110111;
rgb[12296] = 24'b100010001000100010001000;
rgb[12297] = 24'b100110011001100110011001;
rgb[12298] = 24'b101010101010101010101010;
rgb[12299] = 24'b101110111011101110111011;
rgb[12300] = 24'b110011001100110011001100;
rgb[12301] = 24'b110111011101110111011101;
rgb[12302] = 24'b111011101110111011101110;
rgb[12303] = 24'b111111111111111111111111;
rgb[12304] = 24'b000000000000000000000000;
rgb[12305] = 24'b000100010000111100010010;
rgb[12306] = 24'b001000100001111100100100;
rgb[12307] = 24'b001100110010111100110110;
rgb[12308] = 24'b010001000011111101001000;
rgb[12309] = 24'b010101010100111101011010;
rgb[12310] = 24'b011001100101111101101100;
rgb[12311] = 24'b011110000110111101111110;
rgb[12312] = 24'b100010011000000010001111;
rgb[12313] = 24'b100110011001001010011111;
rgb[12314] = 24'b101010101010010010101111;
rgb[12315] = 24'b101110111011011010111111;
rgb[12316] = 24'b110011001100100011001111;
rgb[12317] = 24'b110111011101101011011111;
rgb[12318] = 24'b111011101110110011101111;
rgb[12319] = 24'b111111111111111111111111;
rgb[12320] = 24'b000000000000000000000000;
rgb[12321] = 24'b000100010000111000010011;
rgb[12322] = 24'b001000100001110100100110;
rgb[12323] = 24'b001100110010110000111001;
rgb[12324] = 24'b010001010011101001001101;
rgb[12325] = 24'b010101100100100101100000;
rgb[12326] = 24'b011001110101100001110011;
rgb[12327] = 24'b011110010110011110000110;
rgb[12328] = 24'b100010100111100010010111;
rgb[12329] = 24'b100110101000101110100110;
rgb[12330] = 24'b101010111001111010110101;
rgb[12331] = 24'b101111001011000111000100;
rgb[12332] = 24'b110011001100010111010010;
rgb[12333] = 24'b110111011101100011100001;
rgb[12334] = 24'b111011101110101111110000;
rgb[12335] = 24'b111111111111111111111111;
rgb[12336] = 24'b000000000000000000000000;
rgb[12337] = 24'b000100010000110100010100;
rgb[12338] = 24'b001000100001101100101000;
rgb[12339] = 24'b001101000010100000111101;
rgb[12340] = 24'b010001010011011001010001;
rgb[12341] = 24'b010101110100010001100101;
rgb[12342] = 24'b011010000101000101111010;
rgb[12343] = 24'b011110100101111110001110;
rgb[12344] = 24'b100010110111000010011111;
rgb[12345] = 24'b100110111000010010101101;
rgb[12346] = 24'b101011001001100010111011;
rgb[12347] = 24'b101111001010110111001000;
rgb[12348] = 24'b110011011100000111010110;
rgb[12349] = 24'b110111011101011011100011;
rgb[12350] = 24'b111011101110101011110001;
rgb[12351] = 24'b111111111111111111111111;
rgb[12352] = 24'b000000000000000000000000;
rgb[12353] = 24'b000100010000110000010101;
rgb[12354] = 24'b001000110001100000101011;
rgb[12355] = 24'b001101000010010101000000;
rgb[12356] = 24'b010001100011000101010110;
rgb[12357] = 24'b010110000011111001101011;
rgb[12358] = 24'b011010010100101010000001;
rgb[12359] = 24'b011110110101011110010110;
rgb[12360] = 24'b100011000110100010100111;
rgb[12361] = 24'b100111000111110110110100;
rgb[12362] = 24'b101011011001001111000000;
rgb[12363] = 24'b101111011010100011001101;
rgb[12364] = 24'b110011011011111011011001;
rgb[12365] = 24'b110111101101001111100110;
rgb[12366] = 24'b111011101110100111110010;
rgb[12367] = 24'b111111111111111111111111;
rgb[12368] = 24'b000000000000000000000000;
rgb[12369] = 24'b000100010000101100010110;
rgb[12370] = 24'b001000110001011000101101;
rgb[12371] = 24'b001101010010001001000100;
rgb[12372] = 24'b010001110010110101011010;
rgb[12373] = 24'b010110010011100001110001;
rgb[12374] = 24'b011010100100010010001000;
rgb[12375] = 24'b011111000100111110011110;
rgb[12376] = 24'b100011010110000010101111;
rgb[12377] = 24'b100111010111011010111011;
rgb[12378] = 24'b101011101000110111000110;
rgb[12379] = 24'b101111101010010011010001;
rgb[12380] = 24'b110011101011101111011101;
rgb[12381] = 24'b110111101101000111101000;
rgb[12382] = 24'b111011101110100011110011;
rgb[12383] = 24'b111111111111111111111111;
rgb[12384] = 24'b000000000000000000000000;
rgb[12385] = 24'b000100010000101000010111;
rgb[12386] = 24'b001000110001010000101111;
rgb[12387] = 24'b001101010001111001000111;
rgb[12388] = 24'b010001110010100001011111;
rgb[12389] = 24'b010110010011001101110110;
rgb[12390] = 24'b011010110011110110001110;
rgb[12391] = 24'b011111010100011110100110;
rgb[12392] = 24'b100011100101100010110111;
rgb[12393] = 24'b100111100111000011000001;
rgb[12394] = 24'b101011101000011111001100;
rgb[12395] = 24'b101111101001111111010110;
rgb[12396] = 24'b110011101011011111100000;
rgb[12397] = 24'b110111101100111111101010;
rgb[12398] = 24'b111011101110011111110100;
rgb[12399] = 24'b111111101111111111111110;
rgb[12400] = 24'b000000000000000000000000;
rgb[12401] = 24'b000100100000100100011000;
rgb[12402] = 24'b001001000001001000110001;
rgb[12403] = 24'b001101100001101101001010;
rgb[12404] = 24'b010010000010010001100011;
rgb[12405] = 24'b010110100010110101111100;
rgb[12406] = 24'b011011000011011010010101;
rgb[12407] = 24'b011111100011111110101110;
rgb[12408] = 24'b100011110101000010111111;
rgb[12409] = 24'b100111110110100111001000;
rgb[12410] = 24'b101011111000001011010001;
rgb[12411] = 24'b101111111001101111011010;
rgb[12412] = 24'b110011111011010011100011;
rgb[12413] = 24'b110111111100110111101100;
rgb[12414] = 24'b111011111110011011110101;
rgb[12415] = 24'b111111111111111111111111;
rgb[12416] = 24'b000000000000000000000000;
rgb[12417] = 24'b000100100000011100011010;
rgb[12418] = 24'b001001000000111100110100;
rgb[12419] = 24'b001101100001011101001110;
rgb[12420] = 24'b010010010001111101101000;
rgb[12421] = 24'b010110110010011110000010;
rgb[12422] = 24'b011011010010111110011100;
rgb[12423] = 24'b100000000011011110110110;
rgb[12424] = 24'b100100010100100011000111;
rgb[12425] = 24'b101000000110001011001111;
rgb[12426] = 24'b101100000111110011010111;
rgb[12427] = 24'b110000001001011011011111;
rgb[12428] = 24'b110011111011000011100111;
rgb[12429] = 24'b110111111100101011101111;
rgb[12430] = 24'b111011111110010011110111;
rgb[12431] = 24'b111111101111111111111110;
rgb[12432] = 24'b000000000000000000000000;
rgb[12433] = 24'b000100100000011000011011;
rgb[12434] = 24'b001001000000110100110110;
rgb[12435] = 24'b001101110001010001010001;
rgb[12436] = 24'b010010010001101101101100;
rgb[12437] = 24'b010111000010000110001000;
rgb[12438] = 24'b011011100010100010100011;
rgb[12439] = 24'b100000010010111110111110;
rgb[12440] = 24'b100100100100000011001111;
rgb[12441] = 24'b101000010101101111010110;
rgb[12442] = 24'b101100010111011011011101;
rgb[12443] = 24'b110000001001001011100011;
rgb[12444] = 24'b110100001010110111101010;
rgb[12445] = 24'b110111111100100011110001;
rgb[12446] = 24'b111011111110001111111000;
rgb[12447] = 24'b111111111111111111111111;
rgb[12448] = 24'b000000000000000000000000;
rgb[12449] = 24'b000100100000010100011100;
rgb[12450] = 24'b001001010000101100111000;
rgb[12451] = 24'b001101110001000101010101;
rgb[12452] = 24'b010010100001011001110001;
rgb[12453] = 24'b010111010001110010001101;
rgb[12454] = 24'b011011110010001010101010;
rgb[12455] = 24'b100000100010011111000110;
rgb[12456] = 24'b100100110011100011010111;
rgb[12457] = 24'b101000100101010011011101;
rgb[12458] = 24'b101100100111000111100010;
rgb[12459] = 24'b110000011000110111101000;
rgb[12460] = 24'b110100001010101011101110;
rgb[12461] = 24'b111000001100011011110011;
rgb[12462] = 24'b111011111110001011111001;
rgb[12463] = 24'b111111101111111111111110;
rgb[12464] = 24'b000000000000000000000000;
rgb[12465] = 24'b000100100000010000011101;
rgb[12466] = 24'b001001010000100100111010;
rgb[12467] = 24'b001110000000110101011000;
rgb[12468] = 24'b010010110001001001110101;
rgb[12469] = 24'b010111010001011010010011;
rgb[12470] = 24'b011100000001101110110000;
rgb[12471] = 24'b100000110001111111001110;
rgb[12472] = 24'b100101000011000011011111;
rgb[12473] = 24'b101000110100111011100011;
rgb[12474] = 24'b101100100110101111101000;
rgb[12475] = 24'b110000101000100111101100;
rgb[12476] = 24'b110100011010011011110001;
rgb[12477] = 24'b111000001100010011110101;
rgb[12478] = 24'b111011111110000111111010;
rgb[12479] = 24'b111111111111111111111111;
rgb[12480] = 24'b000000000000000000000000;
rgb[12481] = 24'b000100100000001100011110;
rgb[12482] = 24'b001001010000011000111101;
rgb[12483] = 24'b001110000000101001011011;
rgb[12484] = 24'b010010110000110101111010;
rgb[12485] = 24'b010111100001000010011001;
rgb[12486] = 24'b011100010001010010110111;
rgb[12487] = 24'b100001000001011111010110;
rgb[12488] = 24'b100101010010100011100111;
rgb[12489] = 24'b101001000100011111101010;
rgb[12490] = 24'b101100110110010111101110;
rgb[12491] = 24'b110000101000010011110001;
rgb[12492] = 24'b110100011010001111110100;
rgb[12493] = 24'b111000001100000111111000;
rgb[12494] = 24'b111011111110000011111011;
rgb[12495] = 24'b111111111111111111111111;
rgb[12496] = 24'b000000000000000000000000;
rgb[12497] = 24'b000100110000001000011111;
rgb[12498] = 24'b001001100000010000111111;
rgb[12499] = 24'b001110010000011001011111;
rgb[12500] = 24'b010011000000100101111110;
rgb[12501] = 24'b010111110000101110011110;
rgb[12502] = 24'b011100100000110110111110;
rgb[12503] = 24'b100001010000111111011110;
rgb[12504] = 24'b100101100010000011101111;
rgb[12505] = 24'b101001010100000011110001;
rgb[12506] = 24'b101101000110000011110011;
rgb[12507] = 24'b110000111000000011110101;
rgb[12508] = 24'b110100101001111111111000;
rgb[12509] = 24'b111000011011111111111010;
rgb[12510] = 24'b111100001101111111111100;
rgb[12511] = 24'b111111111111111111111111;
rgb[12512] = 24'b000000000000000000000000;
rgb[12513] = 24'b000100110000000100100000;
rgb[12514] = 24'b001001100000001001000001;
rgb[12515] = 24'b001110010000001101100010;
rgb[12516] = 24'b010011010000010010000011;
rgb[12517] = 24'b011000000000010110100100;
rgb[12518] = 24'b011100110000011011000101;
rgb[12519] = 24'b100001100000011111100110;
rgb[12520] = 24'b100101110001100011110111;
rgb[12521] = 24'b101001100011100111111000;
rgb[12522] = 24'b101101010101101011111001;
rgb[12523] = 24'b110001000111101111111010;
rgb[12524] = 24'b110100101001110011111011;
rgb[12525] = 24'b111000011011110111111100;
rgb[12526] = 24'b111100001101111011111101;
rgb[12527] = 24'b111111111111111111111111;
rgb[12528] = 24'b000000000000000000000000;
rgb[12529] = 24'b000100110000000000100010;
rgb[12530] = 24'b001001100000000001000100;
rgb[12531] = 24'b001110100000000001100110;
rgb[12532] = 24'b010011010000000010001000;
rgb[12533] = 24'b011000010000000010101010;
rgb[12534] = 24'b011101000000000011001100;
rgb[12535] = 24'b100001110000000011101110;
rgb[12536] = 24'b100110000001000111111110;
rgb[12537] = 24'b101001110011001011111111;
rgb[12538] = 24'b101101100101010111111110;
rgb[12539] = 24'b110001000111011011111111;
rgb[12540] = 24'b110100111001100111111111;
rgb[12541] = 24'b111000011011101111111111;
rgb[12542] = 24'b111100001101110111111111;
rgb[12543] = 24'b111111111111111111111111;
rgb[12544] = 24'b000000000000000000000000;
rgb[12545] = 24'b000100010001000100010001;
rgb[12546] = 24'b001000100010001000100010;
rgb[12547] = 24'b001100110011001100110011;
rgb[12548] = 24'b010001000100010001000100;
rgb[12549] = 24'b010101010101010101010101;
rgb[12550] = 24'b011001100110011001100110;
rgb[12551] = 24'b011101110111011101110111;
rgb[12552] = 24'b100010001000100010001000;
rgb[12553] = 24'b100110011001100110011001;
rgb[12554] = 24'b101010101010101010101010;
rgb[12555] = 24'b101110111011101110111011;
rgb[12556] = 24'b110011001100110011001100;
rgb[12557] = 24'b110111011101110111011101;
rgb[12558] = 24'b111011101110111011101110;
rgb[12559] = 24'b111111111111111111111111;
rgb[12560] = 24'b000000000000000000000000;
rgb[12561] = 24'b000100010000111100010010;
rgb[12562] = 24'b001000100001111100100100;
rgb[12563] = 24'b001101000010111100110110;
rgb[12564] = 24'b010001010011111101001000;
rgb[12565] = 24'b010101100100111101011010;
rgb[12566] = 24'b011010000101111101101100;
rgb[12567] = 24'b011110010110111101111110;
rgb[12568] = 24'b100010101000000010001111;
rgb[12569] = 24'b100110111001001010011111;
rgb[12570] = 24'b101010111010010010101111;
rgb[12571] = 24'b101111001011011010111111;
rgb[12572] = 24'b110011011100100011001111;
rgb[12573] = 24'b110111011101101011011111;
rgb[12574] = 24'b111011101110110011101111;
rgb[12575] = 24'b111111111111111111111111;
rgb[12576] = 24'b000000000000000000000000;
rgb[12577] = 24'b000100010000111000010011;
rgb[12578] = 24'b001000110001110100100110;
rgb[12579] = 24'b001101010010110000111001;
rgb[12580] = 24'b010001110011101001001101;
rgb[12581] = 24'b010110000100100101100000;
rgb[12582] = 24'b011010100101100001110011;
rgb[12583] = 24'b011111000110011110000110;
rgb[12584] = 24'b100011010111100010010111;
rgb[12585] = 24'b100111011000101110100110;
rgb[12586] = 24'b101011011001111010110101;
rgb[12587] = 24'b101111101011000111000100;
rgb[12588] = 24'b110011101100010111010010;
rgb[12589] = 24'b110111101101100011100001;
rgb[12590] = 24'b111011101110101111110000;
rgb[12591] = 24'b111111111111111111111111;
rgb[12592] = 24'b000000000000000000000000;
rgb[12593] = 24'b000100100000110100010100;
rgb[12594] = 24'b001001000001101100101000;
rgb[12595] = 24'b001101100010100000111101;
rgb[12596] = 24'b010010000011011001010001;
rgb[12597] = 24'b010110100100010001100101;
rgb[12598] = 24'b011011000101000101111010;
rgb[12599] = 24'b011111100101111110001110;
rgb[12600] = 24'b100011110111000010011111;
rgb[12601] = 24'b100111111000010010101101;
rgb[12602] = 24'b101011111001100010111011;
rgb[12603] = 24'b101111111010110111001000;
rgb[12604] = 24'b110011111100000111010110;
rgb[12605] = 24'b110111111101011011100011;
rgb[12606] = 24'b111011111110101011110001;
rgb[12607] = 24'b111111111111111111111111;
rgb[12608] = 24'b000000000000000000000000;
rgb[12609] = 24'b000100100000110000010101;
rgb[12610] = 24'b001001010001100000101011;
rgb[12611] = 24'b001101110010010101000000;
rgb[12612] = 24'b010010100011000101010110;
rgb[12613] = 24'b010111000011111001101011;
rgb[12614] = 24'b011011110100101010000001;
rgb[12615] = 24'b100000010101011110010110;
rgb[12616] = 24'b100100100110100010100111;
rgb[12617] = 24'b101000100111110110110100;
rgb[12618] = 24'b101100011001001111000000;
rgb[12619] = 24'b110000011010100011001101;
rgb[12620] = 24'b110100001011111011011001;
rgb[12621] = 24'b111000001101001111100110;
rgb[12622] = 24'b111011111110100111110010;
rgb[12623] = 24'b111111111111111111111111;
rgb[12624] = 24'b000000000000000000000000;
rgb[12625] = 24'b000100100000101100010110;
rgb[12626] = 24'b001001010001011000101101;
rgb[12627] = 24'b001110000010001001000100;
rgb[12628] = 24'b010010110010110101011010;
rgb[12629] = 24'b010111100011100001110001;
rgb[12630] = 24'b011100010100010010001000;
rgb[12631] = 24'b100001000100111110011110;
rgb[12632] = 24'b100101010110000010101111;
rgb[12633] = 24'b101001000111011010111011;
rgb[12634] = 24'b101100111000110111000110;
rgb[12635] = 24'b110000101010010011010001;
rgb[12636] = 24'b110100011011101111011101;
rgb[12637] = 24'b111000001101000111101000;
rgb[12638] = 24'b111011111110100011110011;
rgb[12639] = 24'b111111111111111111111111;
rgb[12640] = 24'b000000000000000000000000;
rgb[12641] = 24'b000100110000101000010111;
rgb[12642] = 24'b001001100001010000101111;
rgb[12643] = 24'b001110010001111001000111;
rgb[12644] = 24'b010011010010100001011111;
rgb[12645] = 24'b011000000011001101110110;
rgb[12646] = 24'b011100110011110110001110;
rgb[12647] = 24'b100001100100011110100110;
rgb[12648] = 24'b100101110101100010110111;
rgb[12649] = 24'b101001100111000011000001;
rgb[12650] = 24'b101101011000011111001100;
rgb[12651] = 24'b110001001001111111010110;
rgb[12652] = 24'b110100101011011111100000;
rgb[12653] = 24'b111000011100111111101010;
rgb[12654] = 24'b111100001110011111110100;
rgb[12655] = 24'b111111101111111111111110;
rgb[12656] = 24'b000000000000000000000000;
rgb[12657] = 24'b000100110000100100011000;
rgb[12658] = 24'b001001110001001000110001;
rgb[12659] = 24'b001110100001101101001010;
rgb[12660] = 24'b010011100010010001100011;
rgb[12661] = 24'b011000100010110101111100;
rgb[12662] = 24'b011101010011011010010101;
rgb[12663] = 24'b100010010011111110101110;
rgb[12664] = 24'b100110100101000010111111;
rgb[12665] = 24'b101010000110100111001000;
rgb[12666] = 24'b101101111000001011010001;
rgb[12667] = 24'b110001011001101111011010;
rgb[12668] = 24'b110100111011010011100011;
rgb[12669] = 24'b111000101100110111101100;
rgb[12670] = 24'b111100001110011011110101;
rgb[12671] = 24'b111111111111111111111111;
rgb[12672] = 24'b000000000000000000000000;
rgb[12673] = 24'b000101000000011100011010;
rgb[12674] = 24'b001010000000111100110100;
rgb[12675] = 24'b001111000001011101001110;
rgb[12676] = 24'b010100000001111101101000;
rgb[12677] = 24'b011001000010011110000010;
rgb[12678] = 24'b011110000010111110011100;
rgb[12679] = 24'b100011000011011110110110;
rgb[12680] = 24'b100111010100100011000111;
rgb[12681] = 24'b101010110110001011001111;
rgb[12682] = 24'b101110010111110011010111;
rgb[12683] = 24'b110001111001011011011111;
rgb[12684] = 24'b110101011011000011100111;
rgb[12685] = 24'b111000111100101011101111;
rgb[12686] = 24'b111100011110010011110111;
rgb[12687] = 24'b111111101111111111111110;
rgb[12688] = 24'b000000000000000000000000;
rgb[12689] = 24'b000101000000011000011011;
rgb[12690] = 24'b001010000000110100110110;
rgb[12691] = 24'b001111010001010001010001;
rgb[12692] = 24'b010100010001101101101100;
rgb[12693] = 24'b011001100010000110001000;
rgb[12694] = 24'b011110100010100010100011;
rgb[12695] = 24'b100011100010111110111110;
rgb[12696] = 24'b100111110100000011001111;
rgb[12697] = 24'b101011010101101111010110;
rgb[12698] = 24'b101110110111011011011101;
rgb[12699] = 24'b110010001001001011100011;
rgb[12700] = 24'b110101101010110111101010;
rgb[12701] = 24'b111000111100100011110001;
rgb[12702] = 24'b111100011110001111111000;
rgb[12703] = 24'b111111111111111111111111;
rgb[12704] = 24'b000000000000000000000000;
rgb[12705] = 24'b000101000000010100011100;
rgb[12706] = 24'b001010010000101100111000;
rgb[12707] = 24'b001111100001000101010101;
rgb[12708] = 24'b010100110001011001110001;
rgb[12709] = 24'b011001110001110010001101;
rgb[12710] = 24'b011111000010001010101010;
rgb[12711] = 24'b100100010010011111000110;
rgb[12712] = 24'b101000100011100011010111;
rgb[12713] = 24'b101011110101010011011101;
rgb[12714] = 24'b101111000111000111100010;
rgb[12715] = 24'b110010101000110111101000;
rgb[12716] = 24'b110101111010101011101110;
rgb[12717] = 24'b111001001100011011110011;
rgb[12718] = 24'b111100011110001011111001;
rgb[12719] = 24'b111111101111111111111110;
rgb[12720] = 24'b000000000000000000000000;
rgb[12721] = 24'b000101010000010000011101;
rgb[12722] = 24'b001010100000100100111010;
rgb[12723] = 24'b001111110000110101011000;
rgb[12724] = 24'b010101000001001001110101;
rgb[12725] = 24'b011010010001011010010011;
rgb[12726] = 24'b011111100001101110110000;
rgb[12727] = 24'b100101000001111111001110;
rgb[12728] = 24'b101001010011000011011111;
rgb[12729] = 24'b101100010100111011100011;
rgb[12730] = 24'b101111100110101111101000;
rgb[12731] = 24'b110010111000100111101100;
rgb[12732] = 24'b110110001010011011110001;
rgb[12733] = 24'b111001011100010011110101;
rgb[12734] = 24'b111100101110000111111010;
rgb[12735] = 24'b111111111111111111111111;
rgb[12736] = 24'b000000000000000000000000;
rgb[12737] = 24'b000101010000001100011110;
rgb[12738] = 24'b001010110000011000111101;
rgb[12739] = 24'b010000000000101001011011;
rgb[12740] = 24'b010101100000110101111010;
rgb[12741] = 24'b011010110001000010011001;
rgb[12742] = 24'b100000010001010010110111;
rgb[12743] = 24'b100101100001011111010110;
rgb[12744] = 24'b101001110010100011100111;
rgb[12745] = 24'b101101000100011111101010;
rgb[12746] = 24'b110000000110010111101110;
rgb[12747] = 24'b110011011000010011110001;
rgb[12748] = 24'b110110011010001111110100;
rgb[12749] = 24'b111001101100000111111000;
rgb[12750] = 24'b111100101110000011111011;
rgb[12751] = 24'b111111111111111111111111;
rgb[12752] = 24'b000000000000000000000000;
rgb[12753] = 24'b000101010000001000011111;
rgb[12754] = 24'b001010110000010000111111;
rgb[12755] = 24'b010000010000011001011111;
rgb[12756] = 24'b010101110000100101111110;
rgb[12757] = 24'b011011010000101110011110;
rgb[12758] = 24'b100000110000110110111110;
rgb[12759] = 24'b100110010000111111011110;
rgb[12760] = 24'b101010100010000011101111;
rgb[12761] = 24'b101101100100000011110001;
rgb[12762] = 24'b110000100110000011110011;
rgb[12763] = 24'b110011101000000011110101;
rgb[12764] = 24'b110110101001111111111000;
rgb[12765] = 24'b111001101011111111111010;
rgb[12766] = 24'b111100101101111111111100;
rgb[12767] = 24'b111111111111111111111111;
rgb[12768] = 24'b000000000000000000000000;
rgb[12769] = 24'b000101100000000100100000;
rgb[12770] = 24'b001011000000001001000001;
rgb[12771] = 24'b010000100000001101100010;
rgb[12772] = 24'b010110010000010010000011;
rgb[12773] = 24'b011011110000010110100100;
rgb[12774] = 24'b100001010000011011000101;
rgb[12775] = 24'b100111000000011111100110;
rgb[12776] = 24'b101011010001100011110111;
rgb[12777] = 24'b101110000011100111111000;
rgb[12778] = 24'b110001000101101011111001;
rgb[12779] = 24'b110100000111101111111010;
rgb[12780] = 24'b110110111001110011111011;
rgb[12781] = 24'b111001111011110111111100;
rgb[12782] = 24'b111100111101111011111101;
rgb[12783] = 24'b111111111111111111111111;
rgb[12784] = 24'b000000000000000000000000;
rgb[12785] = 24'b000101100000000000100010;
rgb[12786] = 24'b001011010000000001000100;
rgb[12787] = 24'b010001000000000001100110;
rgb[12788] = 24'b010110100000000010001000;
rgb[12789] = 24'b011100010000000010101010;
rgb[12790] = 24'b100010000000000011001100;
rgb[12791] = 24'b100111100000000011101110;
rgb[12792] = 24'b101011110001000111111110;
rgb[12793] = 24'b101110110011001011111111;
rgb[12794] = 24'b110001100101010111111110;
rgb[12795] = 24'b110100010111011011111111;
rgb[12796] = 24'b110111011001100111111111;
rgb[12797] = 24'b111010001011101111111111;
rgb[12798] = 24'b111100111101110111111111;
rgb[12799] = 24'b111111111111111111111111;
rgb[12800] = 24'b000000000000000000000000;
rgb[12801] = 24'b000100010001000100010001;
rgb[12802] = 24'b001000100010001000100010;
rgb[12803] = 24'b001100110011001100110011;
rgb[12804] = 24'b010001000100010001000100;
rgb[12805] = 24'b010101010101010101010101;
rgb[12806] = 24'b011001100110011001100110;
rgb[12807] = 24'b011101110111011101110111;
rgb[12808] = 24'b100010001000100010001000;
rgb[12809] = 24'b100110011001100110011001;
rgb[12810] = 24'b101010101010101010101010;
rgb[12811] = 24'b101110111011101110111011;
rgb[12812] = 24'b110011001100110011001100;
rgb[12813] = 24'b110111011101110111011101;
rgb[12814] = 24'b111011101110111011101110;
rgb[12815] = 24'b111111111111111111111111;
rgb[12816] = 24'b000000000000000000000000;
rgb[12817] = 24'b000100010000111100010010;
rgb[12818] = 24'b001000110001111100100100;
rgb[12819] = 24'b001101000010111100110110;
rgb[12820] = 24'b010001100011111101001000;
rgb[12821] = 24'b010101110100111101011010;
rgb[12822] = 24'b011010010101111101101100;
rgb[12823] = 24'b011110110110111101111110;
rgb[12824] = 24'b100011001000000010001111;
rgb[12825] = 24'b100111001001001010011111;
rgb[12826] = 24'b101011001010010010101111;
rgb[12827] = 24'b101111011011011010111111;
rgb[12828] = 24'b110011011100100011001111;
rgb[12829] = 24'b110111101101101011011111;
rgb[12830] = 24'b111011101110110011101111;
rgb[12831] = 24'b111111111111111111111111;
rgb[12832] = 24'b000000000000000000000000;
rgb[12833] = 24'b000100100000111000010011;
rgb[12834] = 24'b001001000001110100100110;
rgb[12835] = 24'b001101100010110000111001;
rgb[12836] = 24'b010010000011101001001101;
rgb[12837] = 24'b010110100100100101100000;
rgb[12838] = 24'b011011010101100001110011;
rgb[12839] = 24'b011111110110011110000110;
rgb[12840] = 24'b100100000111100010010111;
rgb[12841] = 24'b101000001000101110100110;
rgb[12842] = 24'b101011111001111010110101;
rgb[12843] = 24'b101111111011000111000100;
rgb[12844] = 24'b110011111100010111010010;
rgb[12845] = 24'b110111111101100011100001;
rgb[12846] = 24'b111011111110101111110000;
rgb[12847] = 24'b111111111111111111111111;
rgb[12848] = 24'b000000000000000000000000;
rgb[12849] = 24'b000100100000110100010100;
rgb[12850] = 24'b001001010001101100101000;
rgb[12851] = 24'b001110000010100000111101;
rgb[12852] = 24'b010010110011011001010001;
rgb[12853] = 24'b010111010100010001100101;
rgb[12854] = 24'b011100000101000101111010;
rgb[12855] = 24'b100000110101111110001110;
rgb[12856] = 24'b100101000111000010011111;
rgb[12857] = 24'b101000111000010010101101;
rgb[12858] = 24'b101100101001100010111011;
rgb[12859] = 24'b110000101010110111001000;
rgb[12860] = 24'b110100011100000111010110;
rgb[12861] = 24'b111000001101011011100011;
rgb[12862] = 24'b111011111110101011110001;
rgb[12863] = 24'b111111111111111111111111;
rgb[12864] = 24'b000000000000000000000000;
rgb[12865] = 24'b000100110000110000010101;
rgb[12866] = 24'b001001100001100000101011;
rgb[12867] = 24'b001110100010010101000000;
rgb[12868] = 24'b010011010011000101010110;
rgb[12869] = 24'b011000000011111001101011;
rgb[12870] = 24'b011101000100101010000001;
rgb[12871] = 24'b100001110101011110010110;
rgb[12872] = 24'b100110000110100010100111;
rgb[12873] = 24'b101001110111110110110100;
rgb[12874] = 24'b101101011001001111000000;
rgb[12875] = 24'b110001001010100011001101;
rgb[12876] = 24'b110100111011111011011001;
rgb[12877] = 24'b111000011101001111100110;
rgb[12878] = 24'b111100001110100111110010;
rgb[12879] = 24'b111111111111111111111111;
rgb[12880] = 24'b000000000000000000000000;
rgb[12881] = 24'b000100110000101100010110;
rgb[12882] = 24'b001001110001011000101101;
rgb[12883] = 24'b001110110010001001000100;
rgb[12884] = 24'b010011110010110101011010;
rgb[12885] = 24'b011000110011100001110001;
rgb[12886] = 24'b011101110100010010001000;
rgb[12887] = 24'b100010110100111110011110;
rgb[12888] = 24'b100111000110000010101111;
rgb[12889] = 24'b101010100111011010111011;
rgb[12890] = 24'b101110001000110111000110;
rgb[12891] = 24'b110001101010010011010001;
rgb[12892] = 24'b110101001011101111011101;
rgb[12893] = 24'b111000101101000111101000;
rgb[12894] = 24'b111100001110100011110011;
rgb[12895] = 24'b111111111111111111111111;
rgb[12896] = 24'b000000000000000000000000;
rgb[12897] = 24'b000101000000101000010111;
rgb[12898] = 24'b001010010001010000101111;
rgb[12899] = 24'b001111010001111001000111;
rgb[12900] = 24'b010100100010100001011111;
rgb[12901] = 24'b011001100011001101110110;
rgb[12902] = 24'b011110110011110110001110;
rgb[12903] = 24'b100011110100011110100110;
rgb[12904] = 24'b101000000101100010110111;
rgb[12905] = 24'b101011100111000011000001;
rgb[12906] = 24'b101110111000011111001100;
rgb[12907] = 24'b110010011001111111010110;
rgb[12908] = 24'b110101101011011111100000;
rgb[12909] = 24'b111001001100111111101010;
rgb[12910] = 24'b111100011110011111110100;
rgb[12911] = 24'b111111101111111111111110;
rgb[12912] = 24'b000000000000000000000000;
rgb[12913] = 24'b000101010000100100011000;
rgb[12914] = 24'b001010100001001000110001;
rgb[12915] = 24'b001111110001101101001010;
rgb[12916] = 24'b010101000010010001100011;
rgb[12917] = 24'b011010010010110101111100;
rgb[12918] = 24'b011111100011011010010101;
rgb[12919] = 24'b100101000011111110101110;
rgb[12920] = 24'b101001010101000010111111;
rgb[12921] = 24'b101100010110100111001000;
rgb[12922] = 24'b101111101000001011010001;
rgb[12923] = 24'b110010111001101111011010;
rgb[12924] = 24'b110110001011010011100011;
rgb[12925] = 24'b111001011100110111101100;
rgb[12926] = 24'b111100101110011011110101;
rgb[12927] = 24'b111111111111111111111111;
rgb[12928] = 24'b000000000000000000000000;
rgb[12929] = 24'b000101010000011100011010;
rgb[12930] = 24'b001010110000111100110100;
rgb[12931] = 24'b010000010001011101001110;
rgb[12932] = 24'b010101100001111101101000;
rgb[12933] = 24'b011011000010011110000010;
rgb[12934] = 24'b100000100010111110011100;
rgb[12935] = 24'b100110000011011110110110;
rgb[12936] = 24'b101010010100100011000111;
rgb[12937] = 24'b101101010110001011001111;
rgb[12938] = 24'b110000010111110011010111;
rgb[12939] = 24'b110011011001011011011111;
rgb[12940] = 24'b110110101011000011100111;
rgb[12941] = 24'b111001101100101011101111;
rgb[12942] = 24'b111100101110010011110111;
rgb[12943] = 24'b111111101111111111111110;
rgb[12944] = 24'b000000000000000000000000;
rgb[12945] = 24'b000101100000011000011011;
rgb[12946] = 24'b001011000000110100110110;
rgb[12947] = 24'b010000110001010001010001;
rgb[12948] = 24'b010110010001101101101100;
rgb[12949] = 24'b011011110010000110001000;
rgb[12950] = 24'b100001100010100010100011;
rgb[12951] = 24'b100111000010111110111110;
rgb[12952] = 24'b101011010100000011001111;
rgb[12953] = 24'b101110010101101111010110;
rgb[12954] = 24'b110001000111011011011101;
rgb[12955] = 24'b110100001001001011100011;
rgb[12956] = 24'b110111001010110111101010;
rgb[12957] = 24'b111001111100100011110001;
rgb[12958] = 24'b111100111110001111111000;
rgb[12959] = 24'b111111111111111111111111;
rgb[12960] = 24'b000000000000000000000000;
rgb[12961] = 24'b000101100000010100011100;
rgb[12962] = 24'b001011010000101100111000;
rgb[12963] = 24'b010001000001000101010101;
rgb[12964] = 24'b010110110001011001110001;
rgb[12965] = 24'b011100100001110010001101;
rgb[12966] = 24'b100010010010001010101010;
rgb[12967] = 24'b101000000010011111000110;
rgb[12968] = 24'b101100010011100011010111;
rgb[12969] = 24'b101111000101010011011101;
rgb[12970] = 24'b110001110111000111100010;
rgb[12971] = 24'b110100101000110111101000;
rgb[12972] = 24'b110111011010101011101110;
rgb[12973] = 24'b111010001100011011110011;
rgb[12974] = 24'b111100111110001011111001;
rgb[12975] = 24'b111111101111111111111110;
rgb[12976] = 24'b000000000000000000000000;
rgb[12977] = 24'b000101110000010000011101;
rgb[12978] = 24'b001011110000100100111010;
rgb[12979] = 24'b010001100000110101011000;
rgb[12980] = 24'b010111100001001001110101;
rgb[12981] = 24'b011101010001011010010011;
rgb[12982] = 24'b100011010001101110110000;
rgb[12983] = 24'b101001000001111111001110;
rgb[12984] = 24'b101101010011000011011111;
rgb[12985] = 24'b110000000100111011100011;
rgb[12986] = 24'b110010100110101111101000;
rgb[12987] = 24'b110101011000100111101100;
rgb[12988] = 24'b110111111010011011110001;
rgb[12989] = 24'b111010101100010011110101;
rgb[12990] = 24'b111101001110000111111010;
rgb[12991] = 24'b111111111111111111111111;
rgb[12992] = 24'b000000000000000000000000;
rgb[12993] = 24'b000110000000001100011110;
rgb[12994] = 24'b001100000000011000111101;
rgb[12995] = 24'b010010000000101001011011;
rgb[12996] = 24'b011000000000110101111010;
rgb[12997] = 24'b011110000001000010011001;
rgb[12998] = 24'b100100000001010010110111;
rgb[12999] = 24'b101010000001011111010110;
rgb[13000] = 24'b101110010010100011100111;
rgb[13001] = 24'b110000110100011111101010;
rgb[13002] = 24'b110011010110010111101110;
rgb[13003] = 24'b110101111000010011110001;
rgb[13004] = 24'b111000011010001111110100;
rgb[13005] = 24'b111010111100000111111000;
rgb[13006] = 24'b111101011110000011111011;
rgb[13007] = 24'b111111111111111111111111;
rgb[13008] = 24'b000000000000000000000000;
rgb[13009] = 24'b000110000000001000011111;
rgb[13010] = 24'b001100010000010000111111;
rgb[13011] = 24'b010010100000011001011111;
rgb[13012] = 24'b011000100000100101111110;
rgb[13013] = 24'b011110110000101110011110;
rgb[13014] = 24'b100101000000110110111110;
rgb[13015] = 24'b101011010000111111011110;
rgb[13016] = 24'b101111100010000011101111;
rgb[13017] = 24'b110001110100000011110001;
rgb[13018] = 24'b110100000110000011110011;
rgb[13019] = 24'b110110011000000011110101;
rgb[13020] = 24'b111000111001111111111000;
rgb[13021] = 24'b111011001011111111111010;
rgb[13022] = 24'b111101011101111111111100;
rgb[13023] = 24'b111111111111111111111111;
rgb[13024] = 24'b000000000000000000000000;
rgb[13025] = 24'b000110010000000100100000;
rgb[13026] = 24'b001100100000001001000001;
rgb[13027] = 24'b010010110000001101100010;
rgb[13028] = 24'b011001010000010010000011;
rgb[13029] = 24'b011111100000010110100100;
rgb[13030] = 24'b100101110000011011000101;
rgb[13031] = 24'b101100010000011111100110;
rgb[13032] = 24'b110000100001100011110111;
rgb[13033] = 24'b110010100011100111111000;
rgb[13034] = 24'b110100110101101011111001;
rgb[13035] = 24'b110111000111101111111010;
rgb[13036] = 24'b111001001001110011111011;
rgb[13037] = 24'b111011011011110111111100;
rgb[13038] = 24'b111101101101111011111101;
rgb[13039] = 24'b111111111111111111111111;
rgb[13040] = 24'b000000000000000000000000;
rgb[13041] = 24'b000110010000000000100010;
rgb[13042] = 24'b001100110000000001000100;
rgb[13043] = 24'b010011010000000001100110;
rgb[13044] = 24'b011001110000000010001000;
rgb[13045] = 24'b100000010000000010101010;
rgb[13046] = 24'b100110110000000011001100;
rgb[13047] = 24'b101101010000000011101110;
rgb[13048] = 24'b110001100001000111111110;
rgb[13049] = 24'b110011100011001011111111;
rgb[13050] = 24'b110101100101010111111110;
rgb[13051] = 24'b110111100111011011111111;
rgb[13052] = 24'b111001101001100111111111;
rgb[13053] = 24'b111011101011101111111111;
rgb[13054] = 24'b111101101101110111111111;
rgb[13055] = 24'b111111111111111111111111;
rgb[13056] = 24'b000000000000000000000000;
rgb[13057] = 24'b000100010001000100010001;
rgb[13058] = 24'b001000100010001000100010;
rgb[13059] = 24'b001100110011001100110011;
rgb[13060] = 24'b010001000100010001000100;
rgb[13061] = 24'b010101010101010101010101;
rgb[13062] = 24'b011001100110011001100110;
rgb[13063] = 24'b011101110111011101110111;
rgb[13064] = 24'b100010001000100010001000;
rgb[13065] = 24'b100110011001100110011001;
rgb[13066] = 24'b101010101010101010101010;
rgb[13067] = 24'b101110111011101110111011;
rgb[13068] = 24'b110011001100110011001100;
rgb[13069] = 24'b110111011101110111011101;
rgb[13070] = 24'b111011101110111011101110;
rgb[13071] = 24'b111111111111111111111111;
rgb[13072] = 24'b000000000000000000000000;
rgb[13073] = 24'b000100010000111100010010;
rgb[13074] = 24'b001000110001111100100100;
rgb[13075] = 24'b001101010010111100110110;
rgb[13076] = 24'b010001110011111101001000;
rgb[13077] = 24'b010110010100111101011010;
rgb[13078] = 24'b011010100101111101101100;
rgb[13079] = 24'b011111000110111101111110;
rgb[13080] = 24'b100011011000000010001111;
rgb[13081] = 24'b100111011001001010011111;
rgb[13082] = 24'b101011101010010010101111;
rgb[13083] = 24'b101111101011011010111111;
rgb[13084] = 24'b110011101100100011001111;
rgb[13085] = 24'b110111101101101011011111;
rgb[13086] = 24'b111011101110110011101111;
rgb[13087] = 24'b111111111111111111111111;
rgb[13088] = 24'b000000000000000000000000;
rgb[13089] = 24'b000100100000111000010011;
rgb[13090] = 24'b001001010001110100100110;
rgb[13091] = 24'b001101110010110000111001;
rgb[13092] = 24'b010010100011101001001101;
rgb[13093] = 24'b010111010100100101100000;
rgb[13094] = 24'b011011110101100001110011;
rgb[13095] = 24'b100000100110011110000110;
rgb[13096] = 24'b100100110111100010010111;
rgb[13097] = 24'b101000101000101110100110;
rgb[13098] = 24'b101100101001111010110101;
rgb[13099] = 24'b110000011011000111000100;
rgb[13100] = 24'b110100001100010111010010;
rgb[13101] = 24'b111000001101100011100001;
rgb[13102] = 24'b111011111110101111110000;
rgb[13103] = 24'b111111111111111111111111;
rgb[13104] = 24'b000000000000000000000000;
rgb[13105] = 24'b000100110000110100010100;
rgb[13106] = 24'b001001100001101100101000;
rgb[13107] = 24'b001110100010100000111101;
rgb[13108] = 24'b010011010011011001010001;
rgb[13109] = 24'b011000010100010001100101;
rgb[13110] = 24'b011101000101000101111010;
rgb[13111] = 24'b100001110101111110001110;
rgb[13112] = 24'b100110010111000010011111;
rgb[13113] = 24'b101001111000010010101101;
rgb[13114] = 24'b101101101001100010111011;
rgb[13115] = 24'b110001001010110111001000;
rgb[13116] = 24'b110100111100000111010110;
rgb[13117] = 24'b111000011101011011100011;
rgb[13118] = 24'b111100001110101011110001;
rgb[13119] = 24'b111111111111111111111111;
rgb[13120] = 24'b000000000000000000000000;
rgb[13121] = 24'b000101000000110000010101;
rgb[13122] = 24'b001010000001100000101011;
rgb[13123] = 24'b001111000010010101000000;
rgb[13124] = 24'b010100000011000101010110;
rgb[13125] = 24'b011001010011111001101011;
rgb[13126] = 24'b011110010100101010000001;
rgb[13127] = 24'b100011010101011110010110;
rgb[13128] = 24'b100111100110100010100111;
rgb[13129] = 24'b101011000111110110110100;
rgb[13130] = 24'b101110101001001111000000;
rgb[13131] = 24'b110001111010100011001101;
rgb[13132] = 24'b110101011011111011011001;
rgb[13133] = 24'b111000111101001111100110;
rgb[13134] = 24'b111100011110100111110010;
rgb[13135] = 24'b111111111111111111111111;
rgb[13136] = 24'b000000000000000000000000;
rgb[13137] = 24'b000101010000101100010110;
rgb[13138] = 24'b001010100001011000101101;
rgb[13139] = 24'b001111110010001001000100;
rgb[13140] = 24'b010101000010110101011010;
rgb[13141] = 24'b011010010011100001110001;
rgb[13142] = 24'b011111100100010010001000;
rgb[13143] = 24'b100100110100111110011110;
rgb[13144] = 24'b101001000110000010101111;
rgb[13145] = 24'b101100010111011010111011;
rgb[13146] = 24'b101111101000110111000110;
rgb[13147] = 24'b110010111010010011010001;
rgb[13148] = 24'b110110001011101111011101;
rgb[13149] = 24'b111001011101000111101000;
rgb[13150] = 24'b111100101110100011110011;
rgb[13151] = 24'b111111111111111111111111;
rgb[13152] = 24'b000000000000000000000000;
rgb[13153] = 24'b000101010000101000010111;
rgb[13154] = 24'b001010110001010000101111;
rgb[13155] = 24'b010000010001111001000111;
rgb[13156] = 24'b010101110010100001011111;
rgb[13157] = 24'b011011010011001101110110;
rgb[13158] = 24'b100000110011110110001110;
rgb[13159] = 24'b100110000100011110100110;
rgb[13160] = 24'b101010010101100010110111;
rgb[13161] = 24'b101101100111000011000001;
rgb[13162] = 24'b110000101000011111001100;
rgb[13163] = 24'b110011101001111111010110;
rgb[13164] = 24'b110110101011011111100000;
rgb[13165] = 24'b111001101100111111101010;
rgb[13166] = 24'b111100101110011111110100;
rgb[13167] = 24'b111111101111111111111110;
rgb[13168] = 24'b000000000000000000000000;
rgb[13169] = 24'b000101100000100100011000;
rgb[13170] = 24'b001011010001001000110001;
rgb[13171] = 24'b010000110001101101001010;
rgb[13172] = 24'b010110100010010001100011;
rgb[13173] = 24'b011100010010110101111100;
rgb[13174] = 24'b100001110011011010010101;
rgb[13175] = 24'b100111100011111110101110;
rgb[13176] = 24'b101011110101000010111111;
rgb[13177] = 24'b101110100110100111001000;
rgb[13178] = 24'b110001101000001011010001;
rgb[13179] = 24'b110100011001101111011010;
rgb[13180] = 24'b110111001011010011100011;
rgb[13181] = 24'b111010001100110111101100;
rgb[13182] = 24'b111100111110011011110101;
rgb[13183] = 24'b111111111111111111111111;
rgb[13184] = 24'b000000000000000000000000;
rgb[13185] = 24'b000101110000011100011010;
rgb[13186] = 24'b001011100000111100110100;
rgb[13187] = 24'b010001100001011101001110;
rgb[13188] = 24'b010111010001111101101000;
rgb[13189] = 24'b011101010010011110000010;
rgb[13190] = 24'b100011000010111110011100;
rgb[13191] = 24'b101001000011011110110110;
rgb[13192] = 24'b101101010100100011000111;
rgb[13193] = 24'b101111110110001011001111;
rgb[13194] = 24'b110010100111110011010111;
rgb[13195] = 24'b110101001001011011011111;
rgb[13196] = 24'b110111111011000011100111;
rgb[13197] = 24'b111010011100101011101111;
rgb[13198] = 24'b111101001110010011110111;
rgb[13199] = 24'b111111101111111111111110;
rgb[13200] = 24'b000000000000000000000000;
rgb[13201] = 24'b000110000000011000011011;
rgb[13202] = 24'b001100000000110100110110;
rgb[13203] = 24'b010010000001010001010001;
rgb[13204] = 24'b011000010001101101101100;
rgb[13205] = 24'b011110010010000110001000;
rgb[13206] = 24'b100100010010100010100011;
rgb[13207] = 24'b101010010010111110111110;
rgb[13208] = 24'b101110100100000011001111;
rgb[13209] = 24'b110001000101101111010110;
rgb[13210] = 24'b110011100111011011011101;
rgb[13211] = 24'b110110001001001011100011;
rgb[13212] = 24'b111000011010110111101010;
rgb[13213] = 24'b111010111100100011110001;
rgb[13214] = 24'b111101011110001111111000;
rgb[13215] = 24'b111111111111111111111111;
rgb[13216] = 24'b000000000000000000000000;
rgb[13217] = 24'b000110010000010100011100;
rgb[13218] = 24'b001100100000101100111000;
rgb[13219] = 24'b010010110001000101010101;
rgb[13220] = 24'b011001000001011001110001;
rgb[13221] = 24'b011111010001110010001101;
rgb[13222] = 24'b100101100010001010101010;
rgb[13223] = 24'b101011110010011111000110;
rgb[13224] = 24'b110000000011100011010111;
rgb[13225] = 24'b110010010101010011011101;
rgb[13226] = 24'b110100100111000111100010;
rgb[13227] = 24'b110110111000110111101000;
rgb[13228] = 24'b111001001010101011101110;
rgb[13229] = 24'b111011011100011011110011;
rgb[13230] = 24'b111101101110001011111001;
rgb[13231] = 24'b111111101111111111111110;
rgb[13232] = 24'b000000000000000000000000;
rgb[13233] = 24'b000110010000010000011101;
rgb[13234] = 24'b001100110000100100111010;
rgb[13235] = 24'b010011010000110101011000;
rgb[13236] = 24'b011001110001001001110101;
rgb[13237] = 24'b100000010001011010010011;
rgb[13238] = 24'b100110110001101110110000;
rgb[13239] = 24'b101101010001111111001110;
rgb[13240] = 24'b110001100011000011011111;
rgb[13241] = 24'b110011100100111011100011;
rgb[13242] = 24'b110101100110101111101000;
rgb[13243] = 24'b110111101000100111101100;
rgb[13244] = 24'b111001101010011011110001;
rgb[13245] = 24'b111011101100010011110101;
rgb[13246] = 24'b111101101110000111111010;
rgb[13247] = 24'b111111111111111111111111;
rgb[13248] = 24'b000000000000000000000000;
rgb[13249] = 24'b000110100000001100011110;
rgb[13250] = 24'b001101010000011000111101;
rgb[13251] = 24'b010100000000101001011011;
rgb[13252] = 24'b011010100000110101111010;
rgb[13253] = 24'b100001010001000010011001;
rgb[13254] = 24'b101000000001010010110111;
rgb[13255] = 24'b101110100001011111010110;
rgb[13256] = 24'b110010110010100011100111;
rgb[13257] = 24'b110100110100011111101010;
rgb[13258] = 24'b110110100110010111101110;
rgb[13259] = 24'b111000011000010011110001;
rgb[13260] = 24'b111010011010001111110100;
rgb[13261] = 24'b111100001100000111111000;
rgb[13262] = 24'b111101111110000011111011;
rgb[13263] = 24'b111111111111111111111111;
rgb[13264] = 24'b000000000000000000000000;
rgb[13265] = 24'b000110110000001000011111;
rgb[13266] = 24'b001101110000010000111111;
rgb[13267] = 24'b010100100000011001011111;
rgb[13268] = 24'b011011100000100101111110;
rgb[13269] = 24'b100010010000101110011110;
rgb[13270] = 24'b101001010000110110111110;
rgb[13271] = 24'b110000000000111111011110;
rgb[13272] = 24'b110100010010000011101111;
rgb[13273] = 24'b110110000100000011110001;
rgb[13274] = 24'b110111100110000011110011;
rgb[13275] = 24'b111001011000000011110101;
rgb[13276] = 24'b111010111001111111111000;
rgb[13277] = 24'b111100101011111111111010;
rgb[13278] = 24'b111110001101111111111100;
rgb[13279] = 24'b111111111111111111111111;
rgb[13280] = 24'b000000000000000000000000;
rgb[13281] = 24'b000111000000000100100000;
rgb[13282] = 24'b001110000000001001000001;
rgb[13283] = 24'b010101000000001101100010;
rgb[13284] = 24'b011100010000010010000011;
rgb[13285] = 24'b100011010000010110100100;
rgb[13286] = 24'b101010010000011011000101;
rgb[13287] = 24'b110001100000011111100110;
rgb[13288] = 24'b110101110001100011110111;
rgb[13289] = 24'b110111000011100111111000;
rgb[13290] = 24'b111000100101101011111001;
rgb[13291] = 24'b111010000111101111111010;
rgb[13292] = 24'b111011011001110011111011;
rgb[13293] = 24'b111100111011110111111100;
rgb[13294] = 24'b111110011101111011111101;
rgb[13295] = 24'b111111111111111111111111;
rgb[13296] = 24'b000000000000000000000000;
rgb[13297] = 24'b000111010000000000100010;
rgb[13298] = 24'b001110100000000001000100;
rgb[13299] = 24'b010101110000000001100110;
rgb[13300] = 24'b011101000000000010001000;
rgb[13301] = 24'b100100010000000010101010;
rgb[13302] = 24'b101011100000000011001100;
rgb[13303] = 24'b110010110000000011101110;
rgb[13304] = 24'b110111000001000111111110;
rgb[13305] = 24'b111000010011001011111111;
rgb[13306] = 24'b111001100101010111111110;
rgb[13307] = 24'b111010110111011011111111;
rgb[13308] = 24'b111100001001100111111111;
rgb[13309] = 24'b111101011011101111111111;
rgb[13310] = 24'b111110101101110111111111;
rgb[13311] = 24'b111111111111111111111111;
rgb[13312] = 24'b000000000000000000000000;
rgb[13313] = 24'b000100010001000100010001;
rgb[13314] = 24'b001000100010001000100010;
rgb[13315] = 24'b001100110011001100110011;
rgb[13316] = 24'b010001000100010001000100;
rgb[13317] = 24'b010101010101010101010101;
rgb[13318] = 24'b011001100110011001100110;
rgb[13319] = 24'b011101110111011101110111;
rgb[13320] = 24'b100010001000100010001000;
rgb[13321] = 24'b100110011001100110011001;
rgb[13322] = 24'b101010101010101010101010;
rgb[13323] = 24'b101110111011101110111011;
rgb[13324] = 24'b110011001100110011001100;
rgb[13325] = 24'b110111011101110111011101;
rgb[13326] = 24'b111011101110111011101110;
rgb[13327] = 24'b111111111111111111111111;
rgb[13328] = 24'b000000000000000000000000;
rgb[13329] = 24'b000100100000111100010010;
rgb[13330] = 24'b001001000001111100100100;
rgb[13331] = 24'b001101100010111100110110;
rgb[13332] = 24'b010010000011111101001000;
rgb[13333] = 24'b010110100100111101011010;
rgb[13334] = 24'b011011000101111101101100;
rgb[13335] = 24'b011111100110111101111110;
rgb[13336] = 24'b100011111000000010001111;
rgb[13337] = 24'b100111111001001010011111;
rgb[13338] = 24'b101011111010010010101111;
rgb[13339] = 24'b101111111011011010111111;
rgb[13340] = 24'b110011111100100011001111;
rgb[13341] = 24'b110111111101101011011111;
rgb[13342] = 24'b111011111110110011101111;
rgb[13343] = 24'b111111111111111111111111;
rgb[13344] = 24'b000000000000000000000000;
rgb[13345] = 24'b000100110000111000010011;
rgb[13346] = 24'b001001100001110100100110;
rgb[13347] = 24'b001110010010110000111001;
rgb[13348] = 24'b010011000011101001001101;
rgb[13349] = 24'b010111110100100101100000;
rgb[13350] = 24'b011100100101100001110011;
rgb[13351] = 24'b100001010110011110000110;
rgb[13352] = 24'b100101100111100010010111;
rgb[13353] = 24'b101001011000101110100110;
rgb[13354] = 24'b101101001001111010110101;
rgb[13355] = 24'b110000111011000111000100;
rgb[13356] = 24'b110100101100010111010010;
rgb[13357] = 24'b111000011101100011100001;
rgb[13358] = 24'b111100001110101111110000;
rgb[13359] = 24'b111111111111111111111111;
rgb[13360] = 24'b000000000000000000000000;
rgb[13361] = 24'b000101000000110100010100;
rgb[13362] = 24'b001010000001101100101000;
rgb[13363] = 24'b001111000010100000111101;
rgb[13364] = 24'b010100000011011001010001;
rgb[13365] = 24'b011001000100010001100101;
rgb[13366] = 24'b011110000101000101111010;
rgb[13367] = 24'b100011000101111110001110;
rgb[13368] = 24'b100111010111000010011111;
rgb[13369] = 24'b101010111000010010101101;
rgb[13370] = 24'b101110011001100010111011;
rgb[13371] = 24'b110001111010110111001000;
rgb[13372] = 24'b110101011100000111010110;
rgb[13373] = 24'b111000111101011011100011;
rgb[13374] = 24'b111100011110101011110001;
rgb[13375] = 24'b111111111111111111111111;
rgb[13376] = 24'b000000000000000000000000;
rgb[13377] = 24'b000101010000110000010101;
rgb[13378] = 24'b001010100001100000101011;
rgb[13379] = 24'b001111110010010101000000;
rgb[13380] = 24'b010101000011000101010110;
rgb[13381] = 24'b011010010011111001101011;
rgb[13382] = 24'b011111100100101010000001;
rgb[13383] = 24'b100100110101011110010110;
rgb[13384] = 24'b101001000110100010100111;
rgb[13385] = 24'b101100010111110110110100;
rgb[13386] = 24'b101111101001001111000000;
rgb[13387] = 24'b110010111010100011001101;
rgb[13388] = 24'b110110001011111011011001;
rgb[13389] = 24'b111001011101001111100110;
rgb[13390] = 24'b111100101110100111110010;
rgb[13391] = 24'b111111111111111111111111;
rgb[13392] = 24'b000000000000000000000000;
rgb[13393] = 24'b000101100000101100010110;
rgb[13394] = 24'b001011000001011000101101;
rgb[13395] = 24'b010000100010001001000100;
rgb[13396] = 24'b010110000010110101011010;
rgb[13397] = 24'b011011100011100001110001;
rgb[13398] = 24'b100001000100010010001000;
rgb[13399] = 24'b100110100100111110011110;
rgb[13400] = 24'b101010110110000010101111;
rgb[13401] = 24'b101101110111011010111011;
rgb[13402] = 24'b110000111000110111000110;
rgb[13403] = 24'b110011111010010011010001;
rgb[13404] = 24'b110110111011101111011101;
rgb[13405] = 24'b111001111101000111101000;
rgb[13406] = 24'b111100111110100011110011;
rgb[13407] = 24'b111111111111111111111111;
rgb[13408] = 24'b000000000000000000000000;
rgb[13409] = 24'b000101110000101000010111;
rgb[13410] = 24'b001011100001010000101111;
rgb[13411] = 24'b010001010001111001000111;
rgb[13412] = 24'b010111000010100001011111;
rgb[13413] = 24'b011100110011001101110110;
rgb[13414] = 24'b100010100011110110001110;
rgb[13415] = 24'b101000100100011110100110;
rgb[13416] = 24'b101100110101100010110111;
rgb[13417] = 24'b101111010111000011000001;
rgb[13418] = 24'b110010001000011111001100;
rgb[13419] = 24'b110100111001111111010110;
rgb[13420] = 24'b110111101011011111100000;
rgb[13421] = 24'b111010011100111111101010;
rgb[13422] = 24'b111101001110011111110100;
rgb[13423] = 24'b111111101111111111111110;
rgb[13424] = 24'b000000000000000000000000;
rgb[13425] = 24'b000110000000100100011000;
rgb[13426] = 24'b001100000001001000110001;
rgb[13427] = 24'b010010000001101101001010;
rgb[13428] = 24'b011000000010010001100011;
rgb[13429] = 24'b011110000010110101111100;
rgb[13430] = 24'b100100010011011010010101;
rgb[13431] = 24'b101010010011111110101110;
rgb[13432] = 24'b101110100101000010111111;
rgb[13433] = 24'b110001000110100111001000;
rgb[13434] = 24'b110011011000001011010001;
rgb[13435] = 24'b110101111001101111011010;
rgb[13436] = 24'b111000011011010011100011;
rgb[13437] = 24'b111010111100110111101100;
rgb[13438] = 24'b111101011110011011110101;
rgb[13439] = 24'b111111111111111111111111;
rgb[13440] = 24'b000000000000000000000000;
rgb[13441] = 24'b000110010000011100011010;
rgb[13442] = 24'b001100100000111100110100;
rgb[13443] = 24'b010010110001011101001110;
rgb[13444] = 24'b011001000001111101101000;
rgb[13445] = 24'b011111100010011110000010;
rgb[13446] = 24'b100101110010111110011100;
rgb[13447] = 24'b101100000011011110110110;
rgb[13448] = 24'b110000010100100011000111;
rgb[13449] = 24'b110010100110001011001111;
rgb[13450] = 24'b110100110111110011010111;
rgb[13451] = 24'b110110111001011011011111;
rgb[13452] = 24'b111001001011000011100111;
rgb[13453] = 24'b111011011100101011101111;
rgb[13454] = 24'b111101101110010011110111;
rgb[13455] = 24'b111111101111111111111110;
rgb[13456] = 24'b000000000000000000000000;
rgb[13457] = 24'b000110100000011000011011;
rgb[13458] = 24'b001101000000110100110110;
rgb[13459] = 24'b010011100001010001010001;
rgb[13460] = 24'b011010000001101101101100;
rgb[13461] = 24'b100000110010000110001000;
rgb[13462] = 24'b100111010010100010100011;
rgb[13463] = 24'b101101110010111110111110;
rgb[13464] = 24'b110010000100000011001111;
rgb[13465] = 24'b110100000101101111010110;
rgb[13466] = 24'b110110000111011011011101;
rgb[13467] = 24'b110111111001001011100011;
rgb[13468] = 24'b111001111010110111101010;
rgb[13469] = 24'b111011111100100011110001;
rgb[13470] = 24'b111101111110001111111000;
rgb[13471] = 24'b111111111111111111111111;
rgb[13472] = 24'b000000000000000000000000;
rgb[13473] = 24'b000110110000010100011100;
rgb[13474] = 24'b001101100000101100111000;
rgb[13475] = 24'b010100010001000101010101;
rgb[13476] = 24'b011011010001011001110001;
rgb[13477] = 24'b100010000001110010001101;
rgb[13478] = 24'b101000110010001010101010;
rgb[13479] = 24'b101111100010011111000110;
rgb[13480] = 24'b110011110011100011010111;
rgb[13481] = 24'b110101100101010011011101;
rgb[13482] = 24'b110111010111000111100010;
rgb[13483] = 24'b111001001000110111101000;
rgb[13484] = 24'b111010101010101011101110;
rgb[13485] = 24'b111100011100011011110011;
rgb[13486] = 24'b111110001110001011111001;
rgb[13487] = 24'b111111101111111111111110;
rgb[13488] = 24'b000000000000000000000000;
rgb[13489] = 24'b000111000000010000011101;
rgb[13490] = 24'b001110000000100100111010;
rgb[13491] = 24'b010101000000110101011000;
rgb[13492] = 24'b011100010001001001110101;
rgb[13493] = 24'b100011010001011010010011;
rgb[13494] = 24'b101010010001101110110000;
rgb[13495] = 24'b110001010001111111001110;
rgb[13496] = 24'b110101100011000011011111;
rgb[13497] = 24'b110111000100111011100011;
rgb[13498] = 24'b111000100110101111101000;
rgb[13499] = 24'b111010001000100111101100;
rgb[13500] = 24'b111011011010011011110001;
rgb[13501] = 24'b111100111100010011110101;
rgb[13502] = 24'b111110011110000111111010;
rgb[13503] = 24'b111111111111111111111111;
rgb[13504] = 24'b000000000000000000000000;
rgb[13505] = 24'b000111010000001100011110;
rgb[13506] = 24'b001110100000011000111101;
rgb[13507] = 24'b010101110000101001011011;
rgb[13508] = 24'b011101010000110101111010;
rgb[13509] = 24'b100100100001000010011001;
rgb[13510] = 24'b101011110001010010110111;
rgb[13511] = 24'b110011010001011111010110;
rgb[13512] = 24'b110111100010100011100111;
rgb[13513] = 24'b111000100100011111101010;
rgb[13514] = 24'b111001110110010111101110;
rgb[13515] = 24'b111011001000010011110001;
rgb[13516] = 24'b111100001010001111110100;
rgb[13517] = 24'b111101011100000111111000;
rgb[13518] = 24'b111110101110000011111011;
rgb[13519] = 24'b111111111111111111111111;
rgb[13520] = 24'b000000000000000000000000;
rgb[13521] = 24'b000111100000001000011111;
rgb[13522] = 24'b001111000000010000111111;
rgb[13523] = 24'b010110100000011001011111;
rgb[13524] = 24'b011110010000100101111110;
rgb[13525] = 24'b100101110000101110011110;
rgb[13526] = 24'b101101010000110110111110;
rgb[13527] = 24'b110101000000111111011110;
rgb[13528] = 24'b111001010010000011101111;
rgb[13529] = 24'b111010000100000011110001;
rgb[13530] = 24'b111011000110000011110011;
rgb[13531] = 24'b111100001000000011110101;
rgb[13532] = 24'b111100111001111111111000;
rgb[13533] = 24'b111101111011111111111010;
rgb[13534] = 24'b111110111101111111111100;
rgb[13535] = 24'b111111111111111111111111;
rgb[13536] = 24'b000000000000000000000000;
rgb[13537] = 24'b000111110000000100100000;
rgb[13538] = 24'b001111100000001001000001;
rgb[13539] = 24'b010111100000001101100010;
rgb[13540] = 24'b011111010000010010000011;
rgb[13541] = 24'b100111000000010110100100;
rgb[13542] = 24'b101111000000011011000101;
rgb[13543] = 24'b110110110000011111100110;
rgb[13544] = 24'b111011000001100011110111;
rgb[13545] = 24'b111011110011100111111000;
rgb[13546] = 24'b111100010101101011111001;
rgb[13547] = 24'b111101000111101111111010;
rgb[13548] = 24'b111101111001110011111011;
rgb[13549] = 24'b111110011011110111111100;
rgb[13550] = 24'b111111001101111011111101;
rgb[13551] = 24'b111111111111111111111111;
rgb[13552] = 24'b000000000000000000000000;
rgb[13553] = 24'b001000000000000000100010;
rgb[13554] = 24'b010000000000000001000100;
rgb[13555] = 24'b011000010000000001100110;
rgb[13556] = 24'b100000010000000010001000;
rgb[13557] = 24'b101000010000000010101010;
rgb[13558] = 24'b110000100000000011001100;
rgb[13559] = 24'b111000100000000011101110;
rgb[13560] = 24'b111100110001000111111110;
rgb[13561] = 24'b111101010011001011111111;
rgb[13562] = 24'b111101100101010111111110;
rgb[13563] = 24'b111110000111011011111111;
rgb[13564] = 24'b111110101001100111111111;
rgb[13565] = 24'b111110111011101111111111;
rgb[13566] = 24'b111111011101110111111111;
rgb[13567] = 24'b111111111111111111111111;
rgb[13568] = 24'b000000000000000000000000;
rgb[13569] = 24'b000100010001000100010001;
rgb[13570] = 24'b001000100010001000100010;
rgb[13571] = 24'b001100110011001100110011;
rgb[13572] = 24'b010001000100010001000100;
rgb[13573] = 24'b010101010101010101010101;
rgb[13574] = 24'b011001100110011001100110;
rgb[13575] = 24'b011101110111011101110111;
rgb[13576] = 24'b100010001000100010001000;
rgb[13577] = 24'b100110011001100110011001;
rgb[13578] = 24'b101010101010101010101010;
rgb[13579] = 24'b101110111011101110111011;
rgb[13580] = 24'b110011001100110011001100;
rgb[13581] = 24'b110111011101110111011101;
rgb[13582] = 24'b111011101110111011101110;
rgb[13583] = 24'b111111111111111111111111;
rgb[13584] = 24'b000000000000000000000000;
rgb[13585] = 24'b000100100000111100010010;
rgb[13586] = 24'b001001000001111100100100;
rgb[13587] = 24'b001101100010111100110110;
rgb[13588] = 24'b010010000011111101001000;
rgb[13589] = 24'b010110100100111101011010;
rgb[13590] = 24'b011011000101111101101100;
rgb[13591] = 24'b011111100110111101111110;
rgb[13592] = 24'b100011111000000010001111;
rgb[13593] = 24'b100111111001001010011111;
rgb[13594] = 24'b101011111010010010101111;
rgb[13595] = 24'b101111111011011010111111;
rgb[13596] = 24'b110011111100100011001111;
rgb[13597] = 24'b110111111101101011011111;
rgb[13598] = 24'b111011111110110011101111;
rgb[13599] = 24'b111111111111111111111111;
rgb[13600] = 24'b000000000000000000000000;
rgb[13601] = 24'b000100110000111000010011;
rgb[13602] = 24'b001001100001110100100110;
rgb[13603] = 24'b001110010010110000111001;
rgb[13604] = 24'b010011010011101001001100;
rgb[13605] = 24'b011000000100100101011111;
rgb[13606] = 24'b011100110101100001110010;
rgb[13607] = 24'b100001100110011110000101;
rgb[13608] = 24'b100101110111100010010110;
rgb[13609] = 24'b101001101000101110100101;
rgb[13610] = 24'b101101011001111010110100;
rgb[13611] = 24'b110001001011000111000011;
rgb[13612] = 24'b110100101100010111010010;
rgb[13613] = 24'b111000011101100011100001;
rgb[13614] = 24'b111100001110101111110000;
rgb[13615] = 24'b111111111111111111111111;
rgb[13616] = 24'b000000000000000000000000;
rgb[13617] = 24'b000101000000110100010100;
rgb[13618] = 24'b001010000001101100101000;
rgb[13619] = 24'b001111010010100000111100;
rgb[13620] = 24'b010100010011011001010000;
rgb[13621] = 24'b011001010100010001100100;
rgb[13622] = 24'b011110100101000101111000;
rgb[13623] = 24'b100011100101111110001100;
rgb[13624] = 24'b100111110111000010011101;
rgb[13625] = 24'b101011011000010010101011;
rgb[13626] = 24'b101110111001100010111001;
rgb[13627] = 24'b110010001010110111000111;
rgb[13628] = 24'b110101101100000111010101;
rgb[13629] = 24'b111000111101011011100011;
rgb[13630] = 24'b111100011110101011110001;
rgb[13631] = 24'b111111111111111111111111;
rgb[13632] = 24'b000000000000000000000000;
rgb[13633] = 24'b000101010000110000010101;
rgb[13634] = 24'b001010110001100000101010;
rgb[13635] = 24'b010000000010010100111111;
rgb[13636] = 24'b010101100011000101010100;
rgb[13637] = 24'b011010110011111001101001;
rgb[13638] = 24'b100000010100101001111110;
rgb[13639] = 24'b100101100101011110010011;
rgb[13640] = 24'b101001110110100010100100;
rgb[13641] = 24'b101101000111110110110001;
rgb[13642] = 24'b110000001001001110111110;
rgb[13643] = 24'b110011011010100011001011;
rgb[13644] = 24'b110110011011111011011000;
rgb[13645] = 24'b111001101101001111100101;
rgb[13646] = 24'b111100101110100111110010;
rgb[13647] = 24'b111111111111111111111111;
rgb[13648] = 24'b000000000000000000000000;
rgb[13649] = 24'b000101100000101100010110;
rgb[13650] = 24'b001011010001011000101100;
rgb[13651] = 24'b010001000010001001000010;
rgb[13652] = 24'b010110100010110101011000;
rgb[13653] = 24'b011100010011100001101110;
rgb[13654] = 24'b100010000100010010000100;
rgb[13655] = 24'b100111100100111110011010;
rgb[13656] = 24'b101011110110000010101011;
rgb[13657] = 24'b101110110111011010110111;
rgb[13658] = 24'b110001101000110111000011;
rgb[13659] = 24'b110100011010010011001111;
rgb[13660] = 24'b110111011011101111011011;
rgb[13661] = 24'b111010001101000111100111;
rgb[13662] = 24'b111100111110100011110011;
rgb[13663] = 24'b111111111111111111111111;
rgb[13664] = 24'b000000000000000000000000;
rgb[13665] = 24'b000101110000101000010111;
rgb[13666] = 24'b001011110001010000101110;
rgb[13667] = 24'b010001110001111001000101;
rgb[13668] = 24'b010111110010100001011100;
rgb[13669] = 24'b011101100011001101110011;
rgb[13670] = 24'b100011100011110110001010;
rgb[13671] = 24'b101001100100011110100010;
rgb[13672] = 24'b101101110101100010110011;
rgb[13673] = 24'b110000010111000010111101;
rgb[13674] = 24'b110011001000011111001000;
rgb[13675] = 24'b110101101001111111010011;
rgb[13676] = 24'b111000001011011111011110;
rgb[13677] = 24'b111010101100111111101001;
rgb[13678] = 24'b111101001110011111110100;
rgb[13679] = 24'b111111101111111111111110;
rgb[13680] = 24'b000000000000000000000000;
rgb[13681] = 24'b000110000000100100011000;
rgb[13682] = 24'b001100010001001000110000;
rgb[13683] = 24'b010010100001101101001000;
rgb[13684] = 24'b011000110010010001100000;
rgb[13685] = 24'b011111000010110101111000;
rgb[13686] = 24'b100101010011011010010001;
rgb[13687] = 24'b101011100011111110101001;
rgb[13688] = 24'b101111110101000010111010;
rgb[13689] = 24'b110010000110100111000100;
rgb[13690] = 24'b110100011000001011001101;
rgb[13691] = 24'b110110101001101111010111;
rgb[13692] = 24'b111000111011010011100001;
rgb[13693] = 24'b111011001100110111101011;
rgb[13694] = 24'b111101011110011011110101;
rgb[13695] = 24'b111111111111111111111111;
rgb[13696] = 24'b000000000000000000000000;
rgb[13697] = 24'b000110100000011100011001;
rgb[13698] = 24'b001101000000111100110010;
rgb[13699] = 24'b010011100001011101001011;
rgb[13700] = 24'b011010000001111101100100;
rgb[13701] = 24'b100000100010011101111110;
rgb[13702] = 24'b100111000010111110010111;
rgb[13703] = 24'b101101100011011110110000;
rgb[13704] = 24'b110001110100100011000001;
rgb[13705] = 24'b110011110110001011001010;
rgb[13706] = 24'b110101110111110011010011;
rgb[13707] = 24'b110111111001011011011011;
rgb[13708] = 24'b111001111011000011100100;
rgb[13709] = 24'b111011111100101011101101;
rgb[13710] = 24'b111101111110010011110110;
rgb[13711] = 24'b111111101111111111111110;
rgb[13712] = 24'b000000000000000000000000;
rgb[13713] = 24'b000110110000011000011010;
rgb[13714] = 24'b001101100000110100110100;
rgb[13715] = 24'b010100010001010001001110;
rgb[13716] = 24'b011011000001101101101000;
rgb[13717] = 24'b100010000010000110000011;
rgb[13718] = 24'b101000110010100010011101;
rgb[13719] = 24'b101111100010111110110111;
rgb[13720] = 24'b110011110100000011001000;
rgb[13721] = 24'b110101100101101111010000;
rgb[13722] = 24'b110111010111011011011000;
rgb[13723] = 24'b111000111001001011011111;
rgb[13724] = 24'b111010101010110111100111;
rgb[13725] = 24'b111100011100100011101111;
rgb[13726] = 24'b111110001110001111110111;
rgb[13727] = 24'b111111111111111111111111;
rgb[13728] = 24'b000000000000000000000000;
rgb[13729] = 24'b000111000000010100011011;
rgb[13730] = 24'b001110000000101100110110;
rgb[13731] = 24'b010101010001000101010001;
rgb[13732] = 24'b011100010001011001101101;
rgb[13733] = 24'b100011010001110010001000;
rgb[13734] = 24'b101010100010001010100011;
rgb[13735] = 24'b110001100010011110111110;
rgb[13736] = 24'b110101110011100011001111;
rgb[13737] = 24'b110111010101010011010110;
rgb[13738] = 24'b111000100111000111011101;
rgb[13739] = 24'b111010001000110111100100;
rgb[13740] = 24'b111011101010101011101010;
rgb[13741] = 24'b111100111100011011110001;
rgb[13742] = 24'b111110011110001011111000;
rgb[13743] = 24'b111111101111111111111110;
rgb[13744] = 24'b000000000000000000000000;
rgb[13745] = 24'b000111010000010000011100;
rgb[13746] = 24'b001110100000100100111000;
rgb[13747] = 24'b010110000000110101010100;
rgb[13748] = 24'b011101010001001001110001;
rgb[13749] = 24'b100100110001011010001101;
rgb[13750] = 24'b101100000001101110101001;
rgb[13751] = 24'b110011100001111111000101;
rgb[13752] = 24'b110111110011000011010110;
rgb[13753] = 24'b111000110100111011011100;
rgb[13754] = 24'b111010000110101111100010;
rgb[13755] = 24'b111011001000100111101000;
rgb[13756] = 24'b111100011010011011101101;
rgb[13757] = 24'b111101011100010011110011;
rgb[13758] = 24'b111110101110000111111001;
rgb[13759] = 24'b111111111111111111111111;
rgb[13760] = 24'b000000000000000000000000;
rgb[13761] = 24'b000111100000001100011101;
rgb[13762] = 24'b001111010000011000111010;
rgb[13763] = 24'b010110110000101001010111;
rgb[13764] = 24'b011110100000110101110101;
rgb[13765] = 24'b100110010001000010010010;
rgb[13766] = 24'b101101110001010010101111;
rgb[13767] = 24'b110101100001011111001101;
rgb[13768] = 24'b111001110010100011011110;
rgb[13769] = 24'b111010100100011111100010;
rgb[13770] = 24'b111011100110010111100111;
rgb[13771] = 24'b111100011000010011101100;
rgb[13772] = 24'b111101001010001111110000;
rgb[13773] = 24'b111110001100000111110101;
rgb[13774] = 24'b111110111110000011111010;
rgb[13775] = 24'b111111111111111111111111;
rgb[13776] = 24'b000000000000000000000000;
rgb[13777] = 24'b000111110000001000011110;
rgb[13778] = 24'b001111110000010000111100;
rgb[13779] = 24'b010111110000011001011010;
rgb[13780] = 24'b011111100000100101111001;
rgb[13781] = 24'b100111100000101110010111;
rgb[13782] = 24'b101111100000110110110101;
rgb[13783] = 24'b110111100000111111010100;
rgb[13784] = 24'b111011110010000011100101;
rgb[13785] = 24'b111100010100000011101000;
rgb[13786] = 24'b111100110110000011101100;
rgb[13787] = 24'b111101011000000011110000;
rgb[13788] = 24'b111110001001111111110011;
rgb[13789] = 24'b111110101011111111110111;
rgb[13790] = 24'b111111001101111111111011;
rgb[13791] = 24'b111111111111111111111111;
rgb[13792] = 24'b000000000000000000000000;
rgb[13793] = 24'b001000000000000100011111;
rgb[13794] = 24'b010000010000001000111110;
rgb[13795] = 24'b011000100000001101011110;
rgb[13796] = 24'b100000110000010001111101;
rgb[13797] = 24'b101001000000010110011100;
rgb[13798] = 24'b110001010000011010111100;
rgb[13799] = 24'b111001100000011111011011;
rgb[13800] = 24'b111101110001100011101100;
rgb[13801] = 24'b111110000011100111101111;
rgb[13802] = 24'b111110010101101011110001;
rgb[13803] = 24'b111110100111101111110100;
rgb[13804] = 24'b111110111001110011110111;
rgb[13805] = 24'b111111001011110111111001;
rgb[13806] = 24'b111111011101111011111100;
rgb[13807] = 24'b111111111111111111111111;
rgb[13808] = 24'b000000000000000000000000;
rgb[13809] = 24'b001000100000000000100000;
rgb[13810] = 24'b010001000000000001000000;
rgb[13811] = 24'b011001100000000001100001;
rgb[13812] = 24'b100010000000000010000001;
rgb[13813] = 24'b101010100000000010100001;
rgb[13814] = 24'b110011000000000011000010;
rgb[13815] = 24'b111011100000000011100010;
rgb[13816] = 24'b111111100001000111110011;
rgb[13817] = 24'b111111110011001011110101;
rgb[13818] = 24'b111111100101010111110110;
rgb[13819] = 24'b111111110111011011111000;
rgb[13820] = 24'b111111111001100111111010;
rgb[13821] = 24'b111111111011101111111011;
rgb[13822] = 24'b111111111101110111111101;
rgb[13823] = 24'b111111111111111111111111;
rgb[13824] = 24'b000000000000000000000000;
rgb[13825] = 24'b000100010001000100010001;
rgb[13826] = 24'b001000100010001000100010;
rgb[13827] = 24'b001100110011001100110011;
rgb[13828] = 24'b010001000100010001000100;
rgb[13829] = 24'b010101010101010101010101;
rgb[13830] = 24'b011001100110011001100110;
rgb[13831] = 24'b011101110111011101110111;
rgb[13832] = 24'b100010001000100010001000;
rgb[13833] = 24'b100110011001100110011001;
rgb[13834] = 24'b101010101010101010101010;
rgb[13835] = 24'b101110111011101110111011;
rgb[13836] = 24'b110011001100110011001100;
rgb[13837] = 24'b110111011101110111011101;
rgb[13838] = 24'b111011101110111011101110;
rgb[13839] = 24'b111111111111111111111111;
rgb[13840] = 24'b000000000000000000000000;
rgb[13841] = 24'b000100100000111100010001;
rgb[13842] = 24'b001001000001111100100011;
rgb[13843] = 24'b001101100010111100110101;
rgb[13844] = 24'b010010000011111101000111;
rgb[13845] = 24'b010110100100111101011001;
rgb[13846] = 24'b011011000101111101101010;
rgb[13847] = 24'b011111100110111101111100;
rgb[13848] = 24'b100011111000000010001101;
rgb[13849] = 24'b100111111001001010011101;
rgb[13850] = 24'b101011111010010010101110;
rgb[13851] = 24'b101111111011011010111110;
rgb[13852] = 24'b110011111100100011001110;
rgb[13853] = 24'b110111111101101011011110;
rgb[13854] = 24'b111011111110110011101110;
rgb[13855] = 24'b111111111111111111111111;
rgb[13856] = 24'b000000000000000000000000;
rgb[13857] = 24'b000100110000111000010010;
rgb[13858] = 24'b001001100001110100100101;
rgb[13859] = 24'b001110010010110000110111;
rgb[13860] = 24'b010011010011101001001010;
rgb[13861] = 24'b011000000100100101011101;
rgb[13862] = 24'b011100110101100001101111;
rgb[13863] = 24'b100001100110011110000010;
rgb[13864] = 24'b100101110111100010010011;
rgb[13865] = 24'b101001101000101110100010;
rgb[13866] = 24'b101101011001111010110010;
rgb[13867] = 24'b110001001011000111000001;
rgb[13868] = 24'b110100101100010111010000;
rgb[13869] = 24'b111000011101100011100000;
rgb[13870] = 24'b111100001110101111101111;
rgb[13871] = 24'b111111111111111111111111;
rgb[13872] = 24'b000000000000000000000000;
rgb[13873] = 24'b000101000000110100010011;
rgb[13874] = 24'b001010000001101100100110;
rgb[13875] = 24'b001111010010100000111010;
rgb[13876] = 24'b010100010011011001001101;
rgb[13877] = 24'b011001010100010001100001;
rgb[13878] = 24'b011110100101000101110100;
rgb[13879] = 24'b100011100101111110001000;
rgb[13880] = 24'b100111110111000010011001;
rgb[13881] = 24'b101011011000010010100111;
rgb[13882] = 24'b101110111001100010110110;
rgb[13883] = 24'b110010001010110111000100;
rgb[13884] = 24'b110101101100000111010011;
rgb[13885] = 24'b111000111101011011100001;
rgb[13886] = 24'b111100011110101011110000;
rgb[13887] = 24'b111111111111111111111111;
rgb[13888] = 24'b000000000000000000000000;
rgb[13889] = 24'b000101010000110000010100;
rgb[13890] = 24'b001010110001100000101000;
rgb[13891] = 24'b010000000010010100111100;
rgb[13892] = 24'b010101100011000101010000;
rgb[13893] = 24'b011010110011111001100101;
rgb[13894] = 24'b100000010100101001111001;
rgb[13895] = 24'b100101100101011110001101;
rgb[13896] = 24'b101001110110100010011110;
rgb[13897] = 24'b101101000111110110101100;
rgb[13898] = 24'b110000001001001110111010;
rgb[13899] = 24'b110011011010100011000111;
rgb[13900] = 24'b110110011011111011010101;
rgb[13901] = 24'b111001101101001111100011;
rgb[13902] = 24'b111100101110100111110001;
rgb[13903] = 24'b111111111111111111111111;
rgb[13904] = 24'b000000000000000000000000;
rgb[13905] = 24'b000101100000101100010101;
rgb[13906] = 24'b001011010001011000101010;
rgb[13907] = 24'b010001000010001000111111;
rgb[13908] = 24'b010110100010110101010100;
rgb[13909] = 24'b011100010011100001101001;
rgb[13910] = 24'b100010000100010001111110;
rgb[13911] = 24'b100111100100111110010011;
rgb[13912] = 24'b101011110110000010100100;
rgb[13913] = 24'b101110110111011010110001;
rgb[13914] = 24'b110001101000110110111110;
rgb[13915] = 24'b110100011010010011001011;
rgb[13916] = 24'b110111011011101111011000;
rgb[13917] = 24'b111010001101000111100101;
rgb[13918] = 24'b111100111110100011110010;
rgb[13919] = 24'b111111111111111111111111;
rgb[13920] = 24'b000000000000000000000000;
rgb[13921] = 24'b000101110000101000010101;
rgb[13922] = 24'b001011110001010000101011;
rgb[13923] = 24'b010001110001111001000001;
rgb[13924] = 24'b010111110010100001010111;
rgb[13925] = 24'b011101100011001101101101;
rgb[13926] = 24'b100011100011110110000011;
rgb[13927] = 24'b101001100100011110011001;
rgb[13928] = 24'b101101110101100010101010;
rgb[13929] = 24'b110000010111000010110110;
rgb[13930] = 24'b110011001000011111000010;
rgb[13931] = 24'b110101101001111111001110;
rgb[13932] = 24'b111000001011011111011010;
rgb[13933] = 24'b111010101100111111100110;
rgb[13934] = 24'b111101001110011111110010;
rgb[13935] = 24'b111111101111111111111110;
rgb[13936] = 24'b000000000000000000000000;
rgb[13937] = 24'b000110000000100100010110;
rgb[13938] = 24'b001100010001001000101101;
rgb[13939] = 24'b010010100001101101000100;
rgb[13940] = 24'b011000110010010001011010;
rgb[13941] = 24'b011111000010110101110001;
rgb[13942] = 24'b100101010011011010001000;
rgb[13943] = 24'b101011100011111110011110;
rgb[13944] = 24'b101111110101000010101111;
rgb[13945] = 24'b110010000110100110111011;
rgb[13946] = 24'b110100011000001011000110;
rgb[13947] = 24'b110110101001101111010001;
rgb[13948] = 24'b111000111011010011011101;
rgb[13949] = 24'b111011001100110111101000;
rgb[13950] = 24'b111101011110011011110011;
rgb[13951] = 24'b111111111111111111111111;
rgb[13952] = 24'b000000000000000000000000;
rgb[13953] = 24'b000110100000011100010111;
rgb[13954] = 24'b001101000000111100101110;
rgb[13955] = 24'b010011100001011101000110;
rgb[13956] = 24'b011010000001111101011101;
rgb[13957] = 24'b100000100010011101110101;
rgb[13958] = 24'b100111000010111110001100;
rgb[13959] = 24'b101101100011011110100100;
rgb[13960] = 24'b110001110100100010110101;
rgb[13961] = 24'b110011110110001010111111;
rgb[13962] = 24'b110101110111110011001010;
rgb[13963] = 24'b110111111001011011010100;
rgb[13964] = 24'b111001111011000011011111;
rgb[13965] = 24'b111011111100101011101001;
rgb[13966] = 24'b111101111110010011110100;
rgb[13967] = 24'b111111101111111111111110;
rgb[13968] = 24'b000000000000000000000000;
rgb[13969] = 24'b000110110000011000011000;
rgb[13970] = 24'b001101100000110100110000;
rgb[13971] = 24'b010100010001010001001000;
rgb[13972] = 24'b011011000001101101100001;
rgb[13973] = 24'b100010000010000101111001;
rgb[13974] = 24'b101000110010100010010001;
rgb[13975] = 24'b101111100010111110101010;
rgb[13976] = 24'b110011110100000010111011;
rgb[13977] = 24'b110101100101101111000100;
rgb[13978] = 24'b110111010111011011001110;
rgb[13979] = 24'b111000111001001011011000;
rgb[13980] = 24'b111010101010110111100001;
rgb[13981] = 24'b111100011100100011101011;
rgb[13982] = 24'b111110001110001111110101;
rgb[13983] = 24'b111111111111111111111111;
rgb[13984] = 24'b000000000000000000000000;
rgb[13985] = 24'b000111000000010100011001;
rgb[13986] = 24'b001110000000101100110010;
rgb[13987] = 24'b010101010001000101001011;
rgb[13988] = 24'b011100010001011001100100;
rgb[13989] = 24'b100011010001110001111101;
rgb[13990] = 24'b101010100010001010010110;
rgb[13991] = 24'b110001100010011110101111;
rgb[13992] = 24'b110101110011100011000000;
rgb[13993] = 24'b110111010101010011001001;
rgb[13994] = 24'b111000100111000111010010;
rgb[13995] = 24'b111010001000110111011011;
rgb[13996] = 24'b111011101010101011100100;
rgb[13997] = 24'b111100111100011011101101;
rgb[13998] = 24'b111110011110001011110110;
rgb[13999] = 24'b111111101111111111111110;
rgb[14000] = 24'b000000000000000000000000;
rgb[14001] = 24'b000111010000010000011001;
rgb[14002] = 24'b001110100000100100110011;
rgb[14003] = 24'b010110000000110101001101;
rgb[14004] = 24'b011101010001001001100111;
rgb[14005] = 24'b100100110001011010000001;
rgb[14006] = 24'b101100000001101110011011;
rgb[14007] = 24'b110011100001111110110101;
rgb[14008] = 24'b110111110011000011000110;
rgb[14009] = 24'b111000110100111011001110;
rgb[14010] = 24'b111010000110101111010110;
rgb[14011] = 24'b111011001000100111011110;
rgb[14012] = 24'b111100011010011011100110;
rgb[14013] = 24'b111101011100010011101110;
rgb[14014] = 24'b111110101110000111110110;
rgb[14015] = 24'b111111111111111111111111;
rgb[14016] = 24'b000000000000000000000000;
rgb[14017] = 24'b000111100000001100011010;
rgb[14018] = 24'b001111010000011000110101;
rgb[14019] = 24'b010110110000101001010000;
rgb[14020] = 24'b011110100000110101101010;
rgb[14021] = 24'b100110010001000010000101;
rgb[14022] = 24'b101101110001010010100000;
rgb[14023] = 24'b110101100001011110111011;
rgb[14024] = 24'b111001110010100011001100;
rgb[14025] = 24'b111010100100011111010011;
rgb[14026] = 24'b111011100110010111011010;
rgb[14027] = 24'b111100011000010011100001;
rgb[14028] = 24'b111101001010001111101001;
rgb[14029] = 24'b111110001100000111110000;
rgb[14030] = 24'b111110111110000011110111;
rgb[14031] = 24'b111111111111111111111111;
rgb[14032] = 24'b000000000000000000000000;
rgb[14033] = 24'b000111110000001000011011;
rgb[14034] = 24'b001111110000010000110111;
rgb[14035] = 24'b010111110000011001010010;
rgb[14036] = 24'b011111100000100101101110;
rgb[14037] = 24'b100111100000101110001001;
rgb[14038] = 24'b101111100000110110100101;
rgb[14039] = 24'b110111100000111111000000;
rgb[14040] = 24'b111011110010000011010001;
rgb[14041] = 24'b111100010100000011011000;
rgb[14042] = 24'b111100110110000011011110;
rgb[14043] = 24'b111101011000000011100101;
rgb[14044] = 24'b111110001001111111101011;
rgb[14045] = 24'b111110101011111111110010;
rgb[14046] = 24'b111111001101111111111000;
rgb[14047] = 24'b111111111111111111111111;
rgb[14048] = 24'b000000000000000000000000;
rgb[14049] = 24'b001000000000000100011100;
rgb[14050] = 24'b010000010000001000111000;
rgb[14051] = 24'b011000100000001101010101;
rgb[14052] = 24'b100000110000010001110001;
rgb[14053] = 24'b101001000000010110001101;
rgb[14054] = 24'b110001010000011010101010;
rgb[14055] = 24'b111001100000011111000110;
rgb[14056] = 24'b111101110001100011010111;
rgb[14057] = 24'b111110000011100111011101;
rgb[14058] = 24'b111110010101101011100010;
rgb[14059] = 24'b111110100111101111101000;
rgb[14060] = 24'b111110111001110011101110;
rgb[14061] = 24'b111111001011110111110011;
rgb[14062] = 24'b111111011101111011111001;
rgb[14063] = 24'b111111111111111111111111;
rgb[14064] = 24'b000000000000000000000000;
rgb[14065] = 24'b001000100000000000011101;
rgb[14066] = 24'b010001000000000000111010;
rgb[14067] = 24'b011001100000000001010111;
rgb[14068] = 24'b100010000000000001110100;
rgb[14069] = 24'b101010100000000010010001;
rgb[14070] = 24'b110011000000000010101110;
rgb[14071] = 24'b111011100000000011001100;
rgb[14072] = 24'b111111100001000111011101;
rgb[14073] = 24'b111111110011001011100001;
rgb[14074] = 24'b111111100101010111100110;
rgb[14075] = 24'b111111110111011011101011;
rgb[14076] = 24'b111111111001100111110000;
rgb[14077] = 24'b111111111011101111110101;
rgb[14078] = 24'b111111111101110111111010;
rgb[14079] = 24'b111111111111111111111111;
rgb[14080] = 24'b000000000000000000000000;
rgb[14081] = 24'b000100010001000100010001;
rgb[14082] = 24'b001000100010001000100010;
rgb[14083] = 24'b001100110011001100110011;
rgb[14084] = 24'b010001000100010001000100;
rgb[14085] = 24'b010101010101010101010101;
rgb[14086] = 24'b011001100110011001100110;
rgb[14087] = 24'b011101110111011101110111;
rgb[14088] = 24'b100010001000100010001000;
rgb[14089] = 24'b100110011001100110011001;
rgb[14090] = 24'b101010101010101010101010;
rgb[14091] = 24'b101110111011101110111011;
rgb[14092] = 24'b110011001100110011001100;
rgb[14093] = 24'b110111011101110111011101;
rgb[14094] = 24'b111011101110111011101110;
rgb[14095] = 24'b111111111111111111111111;
rgb[14096] = 24'b000000000000000000000000;
rgb[14097] = 24'b000100100000111100010001;
rgb[14098] = 24'b001001000001111100100011;
rgb[14099] = 24'b001101100010111100110100;
rgb[14100] = 24'b010010000011111101000110;
rgb[14101] = 24'b010110100100111101010111;
rgb[14102] = 24'b011011000101111101101001;
rgb[14103] = 24'b011111100110111101111011;
rgb[14104] = 24'b100011111000000010001100;
rgb[14105] = 24'b100111111001001010011100;
rgb[14106] = 24'b101011111010010010101100;
rgb[14107] = 24'b101111111011011010111101;
rgb[14108] = 24'b110011111100100011001101;
rgb[14109] = 24'b110111111101101011011110;
rgb[14110] = 24'b111011111110110011101110;
rgb[14111] = 24'b111111111111111111111111;
rgb[14112] = 24'b000000000000000000000000;
rgb[14113] = 24'b000100110000111000010010;
rgb[14114] = 24'b001001100001110100100100;
rgb[14115] = 24'b001110010010110000110110;
rgb[14116] = 24'b010011010011101001001000;
rgb[14117] = 24'b011000000100100101011010;
rgb[14118] = 24'b011100110101100001101101;
rgb[14119] = 24'b100001100110011101111111;
rgb[14120] = 24'b100101110111100010010000;
rgb[14121] = 24'b101001101000101110100000;
rgb[14122] = 24'b101101011001111010101111;
rgb[14123] = 24'b110001001011000110111111;
rgb[14124] = 24'b110100101100010111001111;
rgb[14125] = 24'b111000011101100011011111;
rgb[14126] = 24'b111100001110101111101111;
rgb[14127] = 24'b111111111111111111111111;
rgb[14128] = 24'b000000000000000000000000;
rgb[14129] = 24'b000101000000110100010010;
rgb[14130] = 24'b001010000001101100100101;
rgb[14131] = 24'b001111010010100000111000;
rgb[14132] = 24'b010100010011011001001011;
rgb[14133] = 24'b011001010100010001011101;
rgb[14134] = 24'b011110100101000101110000;
rgb[14135] = 24'b100011100101111110000011;
rgb[14136] = 24'b100111110111000010010100;
rgb[14137] = 24'b101011011000010010100011;
rgb[14138] = 24'b101110111001100010110010;
rgb[14139] = 24'b110010001010110111000010;
rgb[14140] = 24'b110101101100000111010001;
rgb[14141] = 24'b111000111101011011100000;
rgb[14142] = 24'b111100011110101011101111;
rgb[14143] = 24'b111111111111111111111111;
rgb[14144] = 24'b000000000000000000000000;
rgb[14145] = 24'b000101010000110000010011;
rgb[14146] = 24'b001010110001100000100110;
rgb[14147] = 24'b010000000010010100111010;
rgb[14148] = 24'b010101100011000101001101;
rgb[14149] = 24'b011010110011111001100000;
rgb[14150] = 24'b100000010100101001110100;
rgb[14151] = 24'b100101100101011110000111;
rgb[14152] = 24'b101001110110100010011000;
rgb[14153] = 24'b101101000111110110100111;
rgb[14154] = 24'b110000001001001110110101;
rgb[14155] = 24'b110011011010100011000100;
rgb[14156] = 24'b110110011011111011010011;
rgb[14157] = 24'b111001101101001111100001;
rgb[14158] = 24'b111100101110100111110000;
rgb[14159] = 24'b111111111111111111111111;
rgb[14160] = 24'b000000000000000000000000;
rgb[14161] = 24'b000101100000101100010011;
rgb[14162] = 24'b001011010001011000100111;
rgb[14163] = 24'b010001000010001000111011;
rgb[14164] = 24'b010110100010110101001111;
rgb[14165] = 24'b011100010011100001100011;
rgb[14166] = 24'b100010000100010001110111;
rgb[14167] = 24'b100111100100111110001011;
rgb[14168] = 24'b101011110110000010011100;
rgb[14169] = 24'b101110110111011010101010;
rgb[14170] = 24'b110001101000110110111000;
rgb[14171] = 24'b110100011010010011000110;
rgb[14172] = 24'b110111011011101111010100;
rgb[14173] = 24'b111010001101000111100010;
rgb[14174] = 24'b111100111110100011110000;
rgb[14175] = 24'b111111111111111111111111;
rgb[14176] = 24'b000000000000000000000000;
rgb[14177] = 24'b000101110000101000010100;
rgb[14178] = 24'b001011110001010000101001;
rgb[14179] = 24'b010001110001111000111101;
rgb[14180] = 24'b010111110010100001010010;
rgb[14181] = 24'b011101100011001101100110;
rgb[14182] = 24'b100011100011110101111011;
rgb[14183] = 24'b101001100100011110001111;
rgb[14184] = 24'b101101110101100010100000;
rgb[14185] = 24'b110000010111000010101110;
rgb[14186] = 24'b110011001000011110111011;
rgb[14187] = 24'b110101101001111111001001;
rgb[14188] = 24'b111000001011011111010110;
rgb[14189] = 24'b111010101100111111100100;
rgb[14190] = 24'b111101001110011111110001;
rgb[14191] = 24'b111111101111111111111110;
rgb[14192] = 24'b000000000000000000000000;
rgb[14193] = 24'b000110000000100100010101;
rgb[14194] = 24'b001100010001001000101010;
rgb[14195] = 24'b010010100001101100111111;
rgb[14196] = 24'b011000110010010001010100;
rgb[14197] = 24'b011111000010110101101001;
rgb[14198] = 24'b100101010011011001111110;
rgb[14199] = 24'b101011100011111110010100;
rgb[14200] = 24'b101111110101000010100101;
rgb[14201] = 24'b110010000110100110110001;
rgb[14202] = 24'b110100011000001010111110;
rgb[14203] = 24'b110110101001101111001011;
rgb[14204] = 24'b111000111011010011011000;
rgb[14205] = 24'b111011001100110111100101;
rgb[14206] = 24'b111101011110011011110010;
rgb[14207] = 24'b111111111111111111111111;
rgb[14208] = 24'b000000000000000000000000;
rgb[14209] = 24'b000110100000011100010101;
rgb[14210] = 24'b001101000000111100101011;
rgb[14211] = 24'b010011100001011101000001;
rgb[14212] = 24'b011010000001111101010110;
rgb[14213] = 24'b100000100010011101101100;
rgb[14214] = 24'b100111000010111110000010;
rgb[14215] = 24'b101101100011011110011000;
rgb[14216] = 24'b110001110100100010101001;
rgb[14217] = 24'b110011110110001010110101;
rgb[14218] = 24'b110101110111110011000001;
rgb[14219] = 24'b110111111001011011001101;
rgb[14220] = 24'b111001111011000011011010;
rgb[14221] = 24'b111011111100101011100110;
rgb[14222] = 24'b111101111110010011110010;
rgb[14223] = 24'b111111101111111111111110;
rgb[14224] = 24'b000000000000000000000000;
rgb[14225] = 24'b000110110000011000010110;
rgb[14226] = 24'b001101100000110100101100;
rgb[14227] = 24'b010100010001010001000011;
rgb[14228] = 24'b011011000001101101011001;
rgb[14229] = 24'b100010000010000101101111;
rgb[14230] = 24'b101000110010100010000110;
rgb[14231] = 24'b101111100010111110011100;
rgb[14232] = 24'b110011110100000010101101;
rgb[14233] = 24'b110101100101101110111001;
rgb[14234] = 24'b110111010111011011000100;
rgb[14235] = 24'b111000111001001011010000;
rgb[14236] = 24'b111010101010110111011100;
rgb[14237] = 24'b111100011100100011100111;
rgb[14238] = 24'b111110001110001111110011;
rgb[14239] = 24'b111111111111111111111111;
rgb[14240] = 24'b000000000000000000000000;
rgb[14241] = 24'b000111000000010100010110;
rgb[14242] = 24'b001110000000101100101101;
rgb[14243] = 24'b010101010001000101000100;
rgb[14244] = 24'b011100010001011001011011;
rgb[14245] = 24'b100011010001110001110010;
rgb[14246] = 24'b101010100010001010001001;
rgb[14247] = 24'b110001100010011110100000;
rgb[14248] = 24'b110101110011100010110001;
rgb[14249] = 24'b110111010101010010111100;
rgb[14250] = 24'b111000100111000111000111;
rgb[14251] = 24'b111010001000110111010010;
rgb[14252] = 24'b111011101010101011011101;
rgb[14253] = 24'b111100111100011011101000;
rgb[14254] = 24'b111110011110001011110011;
rgb[14255] = 24'b111111101111111111111110;
rgb[14256] = 24'b000000000000000000000000;
rgb[14257] = 24'b000111010000010000010111;
rgb[14258] = 24'b001110100000100100101111;
rgb[14259] = 24'b010110000000110101000110;
rgb[14260] = 24'b011101010001001001011110;
rgb[14261] = 24'b100100110001011001110101;
rgb[14262] = 24'b101100000001101110001101;
rgb[14263] = 24'b110011100001111110100100;
rgb[14264] = 24'b110111110011000010110101;
rgb[14265] = 24'b111000110100111011000000;
rgb[14266] = 24'b111010000110101111001010;
rgb[14267] = 24'b111011001000100111010101;
rgb[14268] = 24'b111100011010011011011111;
rgb[14269] = 24'b111101011100010011101010;
rgb[14270] = 24'b111110101110000111110100;
rgb[14271] = 24'b111111111111111111111111;
rgb[14272] = 24'b000000000000000000000000;
rgb[14273] = 24'b000111100000001100011000;
rgb[14274] = 24'b001111010000011000110000;
rgb[14275] = 24'b010110110000101001001000;
rgb[14276] = 24'b011110100000110101100000;
rgb[14277] = 24'b100110010001000001111000;
rgb[14278] = 24'b101101110001010010010000;
rgb[14279] = 24'b110101100001011110101000;
rgb[14280] = 24'b111001110010100010111001;
rgb[14281] = 24'b111010100100011111000011;
rgb[14282] = 24'b111011100110010111001101;
rgb[14283] = 24'b111100011000010011010111;
rgb[14284] = 24'b111101001010001111100001;
rgb[14285] = 24'b111110001100000111101011;
rgb[14286] = 24'b111110111110000011110101;
rgb[14287] = 24'b111111111111111111111111;
rgb[14288] = 24'b000000000000000000000000;
rgb[14289] = 24'b000111110000001000011000;
rgb[14290] = 24'b001111110000010000110001;
rgb[14291] = 24'b010111110000011001001010;
rgb[14292] = 24'b011111100000100101100010;
rgb[14293] = 24'b100111100000101101111011;
rgb[14294] = 24'b101111100000110110010100;
rgb[14295] = 24'b110111100000111110101101;
rgb[14296] = 24'b111011110010000010111110;
rgb[14297] = 24'b111100010100000011000111;
rgb[14298] = 24'b111100110110000011010000;
rgb[14299] = 24'b111101011000000011011001;
rgb[14300] = 24'b111110001001111111100011;
rgb[14301] = 24'b111110101011111111101100;
rgb[14302] = 24'b111111001101111111110101;
rgb[14303] = 24'b111111111111111111111111;
rgb[14304] = 24'b000000000000000000000000;
rgb[14305] = 24'b001000000000000100011001;
rgb[14306] = 24'b010000010000001000110010;
rgb[14307] = 24'b011000100000001101001011;
rgb[14308] = 24'b100000110000010001100101;
rgb[14309] = 24'b101001000000010101111110;
rgb[14310] = 24'b110001010000011010010111;
rgb[14311] = 24'b111001100000011110110001;
rgb[14312] = 24'b111101110001100011000010;
rgb[14313] = 24'b111110000011100111001010;
rgb[14314] = 24'b111110010101101011010011;
rgb[14315] = 24'b111110100111101111011100;
rgb[14316] = 24'b111110111001110011100100;
rgb[14317] = 24'b111111001011110111101101;
rgb[14318] = 24'b111111011101111011110110;
rgb[14319] = 24'b111111111111111111111111;
rgb[14320] = 24'b000000000000000000000000;
rgb[14321] = 24'b001000100000000000011001;
rgb[14322] = 24'b010001000000000000110011;
rgb[14323] = 24'b011001100000000001001101;
rgb[14324] = 24'b100010000000000001100111;
rgb[14325] = 24'b101010100000000010000001;
rgb[14326] = 24'b110011000000000010011011;
rgb[14327] = 24'b111011100000000010110101;
rgb[14328] = 24'b111111100001000111000110;
rgb[14329] = 24'b111111110011001011001110;
rgb[14330] = 24'b111111100101010111010110;
rgb[14331] = 24'b111111110111011011011110;
rgb[14332] = 24'b111111111001100111100110;
rgb[14333] = 24'b111111111011101111101110;
rgb[14334] = 24'b111111111101110111110110;
rgb[14335] = 24'b111111111111111111111111;
rgb[14336] = 24'b000000000000000000000000;
rgb[14337] = 24'b000100010001000100010001;
rgb[14338] = 24'b001000100010001000100010;
rgb[14339] = 24'b001100110011001100110011;
rgb[14340] = 24'b010001000100010001000100;
rgb[14341] = 24'b010101010101010101010101;
rgb[14342] = 24'b011001100110011001100110;
rgb[14343] = 24'b011101110111011101110111;
rgb[14344] = 24'b100010001000100010001000;
rgb[14345] = 24'b100110011001100110011001;
rgb[14346] = 24'b101010101010101010101010;
rgb[14347] = 24'b101110111011101110111011;
rgb[14348] = 24'b110011001100110011001100;
rgb[14349] = 24'b110111011101110111011101;
rgb[14350] = 24'b111011101110111011101110;
rgb[14351] = 24'b111111111111111111111111;
rgb[14352] = 24'b000000000000000000000000;
rgb[14353] = 24'b000100100000111100010001;
rgb[14354] = 24'b001001000001111100100010;
rgb[14355] = 24'b001101100010111100110100;
rgb[14356] = 24'b010010000011111101000101;
rgb[14357] = 24'b010110100100111101010110;
rgb[14358] = 24'b011011000101111101101000;
rgb[14359] = 24'b011111100110111101111001;
rgb[14360] = 24'b100011111000000010001010;
rgb[14361] = 24'b100111111001001010011011;
rgb[14362] = 24'b101011111010010010101011;
rgb[14363] = 24'b101111111011011010111100;
rgb[14364] = 24'b110011111100100011001101;
rgb[14365] = 24'b110111111101101011011101;
rgb[14366] = 24'b111011111110110011101110;
rgb[14367] = 24'b111111111111111111111111;
rgb[14368] = 24'b000000000000000000000000;
rgb[14369] = 24'b000100110000111000010001;
rgb[14370] = 24'b001001100001110100100011;
rgb[14371] = 24'b001110010010110000110101;
rgb[14372] = 24'b010011010011101001000111;
rgb[14373] = 24'b011000000100100101011000;
rgb[14374] = 24'b011100110101100001101010;
rgb[14375] = 24'b100001100110011101111100;
rgb[14376] = 24'b100101110111100010001101;
rgb[14377] = 24'b101001101000101110011101;
rgb[14378] = 24'b101101011001111010101101;
rgb[14379] = 24'b110001001011000110111110;
rgb[14380] = 24'b110100101100010111001110;
rgb[14381] = 24'b111000011101100011011110;
rgb[14382] = 24'b111100001110101111101110;
rgb[14383] = 24'b111111111111111111111111;
rgb[14384] = 24'b000000000000000000000000;
rgb[14385] = 24'b000101000000110100010010;
rgb[14386] = 24'b001010000001101100100100;
rgb[14387] = 24'b001111010010100000110110;
rgb[14388] = 24'b010100010011011001001000;
rgb[14389] = 24'b011001010100010001011010;
rgb[14390] = 24'b011110100101000101101100;
rgb[14391] = 24'b100011100101111101111110;
rgb[14392] = 24'b100111110111000010001111;
rgb[14393] = 24'b101011011000010010011111;
rgb[14394] = 24'b101110111001100010101111;
rgb[14395] = 24'b110010001010110110111111;
rgb[14396] = 24'b110101101100000111001111;
rgb[14397] = 24'b111000111101011011011111;
rgb[14398] = 24'b111100011110101011101111;
rgb[14399] = 24'b111111111111111111111111;
rgb[14400] = 24'b000000000000000000000000;
rgb[14401] = 24'b000101010000110000010010;
rgb[14402] = 24'b001010110001100000100101;
rgb[14403] = 24'b010000000010010100110111;
rgb[14404] = 24'b010101100011000101001010;
rgb[14405] = 24'b011010110011111001011100;
rgb[14406] = 24'b100000010100101001101111;
rgb[14407] = 24'b100101100101011110000001;
rgb[14408] = 24'b101001110110100010010010;
rgb[14409] = 24'b101101000111110110100010;
rgb[14410] = 24'b110000001001001110110001;
rgb[14411] = 24'b110011011010100011000001;
rgb[14412] = 24'b110110011011111011010000;
rgb[14413] = 24'b111001101101001111100000;
rgb[14414] = 24'b111100101110100111101111;
rgb[14415] = 24'b111111111111111111111111;
rgb[14416] = 24'b000000000000000000000000;
rgb[14417] = 24'b000101100000101100010010;
rgb[14418] = 24'b001011010001011000100101;
rgb[14419] = 24'b010001000010001000111000;
rgb[14420] = 24'b010110100010110101001011;
rgb[14421] = 24'b011100010011100001011110;
rgb[14422] = 24'b100010000100010001110001;
rgb[14423] = 24'b100111100100111110000100;
rgb[14424] = 24'b101011110110000010010101;
rgb[14425] = 24'b101110110111011010100100;
rgb[14426] = 24'b110001101000110110110011;
rgb[14427] = 24'b110100011010010011000010;
rgb[14428] = 24'b110111011011101111010001;
rgb[14429] = 24'b111010001101000111100000;
rgb[14430] = 24'b111100111110100011101111;
rgb[14431] = 24'b111111111111111111111111;
rgb[14432] = 24'b000000000000000000000000;
rgb[14433] = 24'b000101110000101000010011;
rgb[14434] = 24'b001011110001010000100110;
rgb[14435] = 24'b010001110001111000111001;
rgb[14436] = 24'b010111110010100001001101;
rgb[14437] = 24'b011101100011001101100000;
rgb[14438] = 24'b100011100011110101110011;
rgb[14439] = 24'b101001100100011110000110;
rgb[14440] = 24'b101101110101100010010111;
rgb[14441] = 24'b110000010111000010100110;
rgb[14442] = 24'b110011001000011110110101;
rgb[14443] = 24'b110101101001111111000100;
rgb[14444] = 24'b111000001011011111010010;
rgb[14445] = 24'b111010101100111111100001;
rgb[14446] = 24'b111101001110011111110000;
rgb[14447] = 24'b111111101111111111111110;
rgb[14448] = 24'b000000000000000000000000;
rgb[14449] = 24'b000110000000100100010011;
rgb[14450] = 24'b001100010001001000100111;
rgb[14451] = 24'b010010100001101100111010;
rgb[14452] = 24'b011000110010010001001110;
rgb[14453] = 24'b011111000010110101100010;
rgb[14454] = 24'b100101010011011001110101;
rgb[14455] = 24'b101011100011111110001001;
rgb[14456] = 24'b101111110101000010011010;
rgb[14457] = 24'b110010000110100110101000;
rgb[14458] = 24'b110100011000001010110111;
rgb[14459] = 24'b110110101001101111000101;
rgb[14460] = 24'b111000111011010011010011;
rgb[14461] = 24'b111011001100110111100010;
rgb[14462] = 24'b111101011110011011110000;
rgb[14463] = 24'b111111111111111111111111;
rgb[14464] = 24'b000000000000000000000000;
rgb[14465] = 24'b000110100000011100010100;
rgb[14466] = 24'b001101000000111100101000;
rgb[14467] = 24'b010011100001011100111100;
rgb[14468] = 24'b011010000001111101010000;
rgb[14469] = 24'b100000100010011101100100;
rgb[14470] = 24'b100111000010111101111000;
rgb[14471] = 24'b101101100011011110001100;
rgb[14472] = 24'b110001110100100010011101;
rgb[14473] = 24'b110011110110001010101011;
rgb[14474] = 24'b110101110111110010111001;
rgb[14475] = 24'b110111111001011011000111;
rgb[14476] = 24'b111001111011000011010101;
rgb[14477] = 24'b111011111100101011100011;
rgb[14478] = 24'b111101111110010011110001;
rgb[14479] = 24'b111111101111111111111110;
rgb[14480] = 24'b000000000000000000000000;
rgb[14481] = 24'b000110110000011000010100;
rgb[14482] = 24'b001101100000110100101000;
rgb[14483] = 24'b010100010001010000111101;
rgb[14484] = 24'b011011000001101101010001;
rgb[14485] = 24'b100010000010000101100101;
rgb[14486] = 24'b101000110010100001111010;
rgb[14487] = 24'b101111100010111110001110;
rgb[14488] = 24'b110011110100000010011111;
rgb[14489] = 24'b110101100101101110101101;
rgb[14490] = 24'b110111010111011010111010;
rgb[14491] = 24'b111000111001001011001000;
rgb[14492] = 24'b111010101010110111010110;
rgb[14493] = 24'b111100011100100011100011;
rgb[14494] = 24'b111110001110001111110001;
rgb[14495] = 24'b111111111111111111111111;
rgb[14496] = 24'b000000000000000000000000;
rgb[14497] = 24'b000111000000010100010100;
rgb[14498] = 24'b001110000000101100101001;
rgb[14499] = 24'b010101010001000100111110;
rgb[14500] = 24'b011100010001011001010011;
rgb[14501] = 24'b100011010001110001100111;
rgb[14502] = 24'b101010100010001001111100;
rgb[14503] = 24'b110001100010011110010001;
rgb[14504] = 24'b110101110011100010100010;
rgb[14505] = 24'b110111010101010010101111;
rgb[14506] = 24'b111000100111000110111100;
rgb[14507] = 24'b111010001000110111001010;
rgb[14508] = 24'b111011101010101011010111;
rgb[14509] = 24'b111100111100011011100100;
rgb[14510] = 24'b111110011110001011110001;
rgb[14511] = 24'b111111101111111111111110;
rgb[14512] = 24'b000000000000000000000000;
rgb[14513] = 24'b000111010000010000010101;
rgb[14514] = 24'b001110100000100100101010;
rgb[14515] = 24'b010110000000110100111111;
rgb[14516] = 24'b011101010001001001010100;
rgb[14517] = 24'b100100110001011001101001;
rgb[14518] = 24'b101100000001101101111110;
rgb[14519] = 24'b110011100001111110010100;
rgb[14520] = 24'b110111110011000010100101;
rgb[14521] = 24'b111000110100111010110001;
rgb[14522] = 24'b111010000110101110111110;
rgb[14523] = 24'b111011001000100111001011;
rgb[14524] = 24'b111100011010011011011000;
rgb[14525] = 24'b111101011100010011100101;
rgb[14526] = 24'b111110101110000111110010;
rgb[14527] = 24'b111111111111111111111111;
rgb[14528] = 24'b000000000000000000000000;
rgb[14529] = 24'b000111100000001100010101;
rgb[14530] = 24'b001111010000011000101011;
rgb[14531] = 24'b010110110000101001000000;
rgb[14532] = 24'b011110100000110101010110;
rgb[14533] = 24'b100110010001000001101011;
rgb[14534] = 24'b101101110001010010000001;
rgb[14535] = 24'b110101100001011110010110;
rgb[14536] = 24'b111001110010100010100111;
rgb[14537] = 24'b111010100100011110110100;
rgb[14538] = 24'b111011100110010111000000;
rgb[14539] = 24'b111100011000010011001101;
rgb[14540] = 24'b111101001010001111011001;
rgb[14541] = 24'b111110001100000111100110;
rgb[14542] = 24'b111110111110000011110010;
rgb[14543] = 24'b111111111111111111111111;
rgb[14544] = 24'b000000000000000000000000;
rgb[14545] = 24'b000111110000001000010101;
rgb[14546] = 24'b001111110000010000101011;
rgb[14547] = 24'b010111110000011001000001;
rgb[14548] = 24'b011111100000100101010111;
rgb[14549] = 24'b100111100000101101101101;
rgb[14550] = 24'b101111100000110110000011;
rgb[14551] = 24'b110111100000111110011001;
rgb[14552] = 24'b111011110010000010101010;
rgb[14553] = 24'b111100010100000010110110;
rgb[14554] = 24'b111100110110000011000010;
rgb[14555] = 24'b111101011000000011001110;
rgb[14556] = 24'b111110001001111111011010;
rgb[14557] = 24'b111110101011111111100110;
rgb[14558] = 24'b111111001101111111110010;
rgb[14559] = 24'b111111111111111111111111;
rgb[14560] = 24'b000000000000000000000000;
rgb[14561] = 24'b001000000000000100010110;
rgb[14562] = 24'b010000010000001000101100;
rgb[14563] = 24'b011000100000001101000010;
rgb[14564] = 24'b100000110000010001011001;
rgb[14565] = 24'b101001000000010101101111;
rgb[14566] = 24'b110001010000011010000101;
rgb[14567] = 24'b111001100000011110011100;
rgb[14568] = 24'b111101110001100010101101;
rgb[14569] = 24'b111110000011100110111000;
rgb[14570] = 24'b111110010101101011000100;
rgb[14571] = 24'b111110100111101111010000;
rgb[14572] = 24'b111110111001110011011011;
rgb[14573] = 24'b111111001011110111100111;
rgb[14574] = 24'b111111011101111011110011;
rgb[14575] = 24'b111111111111111111111111;
rgb[14576] = 24'b000000000000000000000000;
rgb[14577] = 24'b001000100000000000010110;
rgb[14578] = 24'b010001000000000000101101;
rgb[14579] = 24'b011001100000000001000011;
rgb[14580] = 24'b100010000000000001011010;
rgb[14581] = 24'b101010100000000001110001;
rgb[14582] = 24'b110011000000000010000111;
rgb[14583] = 24'b111011100000000010011110;
rgb[14584] = 24'b111111100001000110101111;
rgb[14585] = 24'b111111110011001010111010;
rgb[14586] = 24'b111111100101010111000110;
rgb[14587] = 24'b111111110111011011010001;
rgb[14588] = 24'b111111111001100111011100;
rgb[14589] = 24'b111111111011101111101000;
rgb[14590] = 24'b111111111101110111110011;
rgb[14591] = 24'b111111111111111111111111;
rgb[14592] = 24'b000000000000000000000000;
rgb[14593] = 24'b000100010001000100010001;
rgb[14594] = 24'b001000100010001000100010;
rgb[14595] = 24'b001100110011001100110011;
rgb[14596] = 24'b010001000100010001000100;
rgb[14597] = 24'b010101010101010101010101;
rgb[14598] = 24'b011001100110011001100110;
rgb[14599] = 24'b011101110111011101110111;
rgb[14600] = 24'b100010001000100010001000;
rgb[14601] = 24'b100110011001100110011001;
rgb[14602] = 24'b101010101010101010101010;
rgb[14603] = 24'b101110111011101110111011;
rgb[14604] = 24'b110011001100110011001100;
rgb[14605] = 24'b110111011101110111011101;
rgb[14606] = 24'b111011101110111011101110;
rgb[14607] = 24'b111111111111111111111111;
rgb[14608] = 24'b000000000000000000000000;
rgb[14609] = 24'b000100100000111100010001;
rgb[14610] = 24'b001001000001111100100010;
rgb[14611] = 24'b001101100010111100110011;
rgb[14612] = 24'b010010000011111101000100;
rgb[14613] = 24'b010110100100111101010101;
rgb[14614] = 24'b011011000101111101100110;
rgb[14615] = 24'b011111100110111101111000;
rgb[14616] = 24'b100011111000000010001001;
rgb[14617] = 24'b100111111001001010011001;
rgb[14618] = 24'b101011111010010010101010;
rgb[14619] = 24'b101111111011011010111011;
rgb[14620] = 24'b110011111100100011001100;
rgb[14621] = 24'b110111111101101011011101;
rgb[14622] = 24'b111011111110110011101110;
rgb[14623] = 24'b111111111111111111111111;
rgb[14624] = 24'b000000000000000000000000;
rgb[14625] = 24'b000100110000111000010001;
rgb[14626] = 24'b001001100001110100100010;
rgb[14627] = 24'b001110010010110000110011;
rgb[14628] = 24'b010011010011101001000101;
rgb[14629] = 24'b011000000100100101010110;
rgb[14630] = 24'b011100110101100001100111;
rgb[14631] = 24'b100001100110011101111001;
rgb[14632] = 24'b100101110111100010001010;
rgb[14633] = 24'b101001101000101110011010;
rgb[14634] = 24'b101101011001111010101011;
rgb[14635] = 24'b110001001011000110111100;
rgb[14636] = 24'b110100101100010111001100;
rgb[14637] = 24'b111000011101100011011101;
rgb[14638] = 24'b111100001110101111101110;
rgb[14639] = 24'b111111111111111111111111;
rgb[14640] = 24'b000000000000000000000000;
rgb[14641] = 24'b000101000000110100010001;
rgb[14642] = 24'b001010000001101100100010;
rgb[14643] = 24'b001111010010100000110100;
rgb[14644] = 24'b010100010011011001000101;
rgb[14645] = 24'b011001010100010001010111;
rgb[14646] = 24'b011110100101000101101000;
rgb[14647] = 24'b100011100101111101111010;
rgb[14648] = 24'b100111110111000010001011;
rgb[14649] = 24'b101011011000010010011011;
rgb[14650] = 24'b101110111001100010101100;
rgb[14651] = 24'b110010001010110110111100;
rgb[14652] = 24'b110101101100000111001101;
rgb[14653] = 24'b111000111101011011011101;
rgb[14654] = 24'b111100011110101011101110;
rgb[14655] = 24'b111111111111111111111111;
rgb[14656] = 24'b000000000000000000000000;
rgb[14657] = 24'b000101010000110000010001;
rgb[14658] = 24'b001010110001100000100011;
rgb[14659] = 24'b010000000010010100110100;
rgb[14660] = 24'b010101100011000101000110;
rgb[14661] = 24'b011010110011111001011000;
rgb[14662] = 24'b100000010100101001101001;
rgb[14663] = 24'b100101100101011101111011;
rgb[14664] = 24'b101001110110100010001100;
rgb[14665] = 24'b101101000111110110011100;
rgb[14666] = 24'b110000001001001110101101;
rgb[14667] = 24'b110011011010100010111101;
rgb[14668] = 24'b110110011011111011001101;
rgb[14669] = 24'b111001101101001111011110;
rgb[14670] = 24'b111100101110100111101110;
rgb[14671] = 24'b111111111111111111111111;
rgb[14672] = 24'b000000000000000000000000;
rgb[14673] = 24'b000101100000101100010001;
rgb[14674] = 24'b001011010001011000100011;
rgb[14675] = 24'b010001000010001000110101;
rgb[14676] = 24'b010110100010110101000111;
rgb[14677] = 24'b011100010011100001011001;
rgb[14678] = 24'b100010000100010001101010;
rgb[14679] = 24'b100111100100111101111100;
rgb[14680] = 24'b101011110110000010001101;
rgb[14681] = 24'b101110110111011010011101;
rgb[14682] = 24'b110001101000110110101110;
rgb[14683] = 24'b110100011010010010111110;
rgb[14684] = 24'b110111011011101111001110;
rgb[14685] = 24'b111010001101000111011110;
rgb[14686] = 24'b111100111110100011101110;
rgb[14687] = 24'b111111111111111111111111;
rgb[14688] = 24'b000000000000000000000000;
rgb[14689] = 24'b000101110000101000010001;
rgb[14690] = 24'b001011110001010000100011;
rgb[14691] = 24'b010001110001111000110101;
rgb[14692] = 24'b010111110010100001000111;
rgb[14693] = 24'b011101100011001101011001;
rgb[14694] = 24'b100011100011110101101011;
rgb[14695] = 24'b101001100100011101111101;
rgb[14696] = 24'b101101110101100010001110;
rgb[14697] = 24'b110000010111000010011110;
rgb[14698] = 24'b110011001000011110101110;
rgb[14699] = 24'b110101101001111110111110;
rgb[14700] = 24'b111000001011011111001110;
rgb[14701] = 24'b111010101100111111011110;
rgb[14702] = 24'b111101001110011111101110;
rgb[14703] = 24'b111111101111111111111110;
rgb[14704] = 24'b000000000000000000000000;
rgb[14705] = 24'b000110000000100100010010;
rgb[14706] = 24'b001100010001001000100100;
rgb[14707] = 24'b010010100001101100110110;
rgb[14708] = 24'b011000110010010001001000;
rgb[14709] = 24'b011111000010110101011010;
rgb[14710] = 24'b100101010011011001101100;
rgb[14711] = 24'b101011100011111101111110;
rgb[14712] = 24'b101111110101000010001111;
rgb[14713] = 24'b110010000110100110011111;
rgb[14714] = 24'b110100011000001010101111;
rgb[14715] = 24'b110110101001101110111111;
rgb[14716] = 24'b111000111011010011001111;
rgb[14717] = 24'b111011001100110111011111;
rgb[14718] = 24'b111101011110011011101111;
rgb[14719] = 24'b111111111111111111111111;
rgb[14720] = 24'b000000000000000000000000;
rgb[14721] = 24'b000110100000011100010010;
rgb[14722] = 24'b001101000000111100100100;
rgb[14723] = 24'b010011100001011100110110;
rgb[14724] = 24'b011010000001111101001001;
rgb[14725] = 24'b100000100010011101011011;
rgb[14726] = 24'b100111000010111101101101;
rgb[14727] = 24'b101101100011011110000000;
rgb[14728] = 24'b110001110100100010010001;
rgb[14729] = 24'b110011110110001010100000;
rgb[14730] = 24'b110101110111110010110000;
rgb[14731] = 24'b110111111001011011000000;
rgb[14732] = 24'b111001111011000011001111;
rgb[14733] = 24'b111011111100101011011111;
rgb[14734] = 24'b111101111110010011101111;
rgb[14735] = 24'b111111101111111111111110;
rgb[14736] = 24'b000000000000000000000000;
rgb[14737] = 24'b000110110000011000010010;
rgb[14738] = 24'b001101100000110100100100;
rgb[14739] = 24'b010100010001010000110111;
rgb[14740] = 24'b011011000001101101001001;
rgb[14741] = 24'b100010000010000101011100;
rgb[14742] = 24'b101000110010100001101110;
rgb[14743] = 24'b101111100010111110000001;
rgb[14744] = 24'b110011110100000010010010;
rgb[14745] = 24'b110101100101101110100001;
rgb[14746] = 24'b110111010111011010110001;
rgb[14747] = 24'b111000111001001011000000;
rgb[14748] = 24'b111010101010110111010000;
rgb[14749] = 24'b111100011100100011011111;
rgb[14750] = 24'b111110001110001111101111;
rgb[14751] = 24'b111111111111111111111111;
rgb[14752] = 24'b000000000000000000000000;
rgb[14753] = 24'b000111000000010100010010;
rgb[14754] = 24'b001110000000101100100101;
rgb[14755] = 24'b010101010001000100110111;
rgb[14756] = 24'b011100010001011001001010;
rgb[14757] = 24'b100011010001110001011101;
rgb[14758] = 24'b101010100010001001101111;
rgb[14759] = 24'b110001100010011110000010;
rgb[14760] = 24'b110101110011100010010011;
rgb[14761] = 24'b110111010101010010100010;
rgb[14762] = 24'b111000100111000110110010;
rgb[14763] = 24'b111010001000110111000001;
rgb[14764] = 24'b111011101010101011010000;
rgb[14765] = 24'b111100111100011011100000;
rgb[14766] = 24'b111110011110001011101111;
rgb[14767] = 24'b111111101111111111111110;
rgb[14768] = 24'b000000000000000000000000;
rgb[14769] = 24'b000111010000010000010010;
rgb[14770] = 24'b001110100000100100100101;
rgb[14771] = 24'b010110000000110100111000;
rgb[14772] = 24'b011101010001001001001011;
rgb[14773] = 24'b100100110001011001011101;
rgb[14774] = 24'b101100000001101101110000;
rgb[14775] = 24'b110011100001111110000011;
rgb[14776] = 24'b110111110011000010010100;
rgb[14777] = 24'b111000110100111010100011;
rgb[14778] = 24'b111010000110101110110010;
rgb[14779] = 24'b111011001000100111000010;
rgb[14780] = 24'b111100011010011011010001;
rgb[14781] = 24'b111101011100010011100000;
rgb[14782] = 24'b111110101110000111101111;
rgb[14783] = 24'b111111111111111111111111;
rgb[14784] = 24'b000000000000000000000000;
rgb[14785] = 24'b000111100000001100010010;
rgb[14786] = 24'b001111010000011000100101;
rgb[14787] = 24'b010110110000101000111000;
rgb[14788] = 24'b011110100000110101001011;
rgb[14789] = 24'b100110010001000001011110;
rgb[14790] = 24'b101101110001010001110001;
rgb[14791] = 24'b110101100001011110000100;
rgb[14792] = 24'b111001110010100010010101;
rgb[14793] = 24'b111010100100011110100100;
rgb[14794] = 24'b111011100110010110110011;
rgb[14795] = 24'b111100011000010011000010;
rgb[14796] = 24'b111101001010001111010001;
rgb[14797] = 24'b111110001100000111100000;
rgb[14798] = 24'b111110111110000011101111;
rgb[14799] = 24'b111111111111111111111111;
rgb[14800] = 24'b000000000000000000000000;
rgb[14801] = 24'b000111110000001000010011;
rgb[14802] = 24'b001111110000010000100110;
rgb[14803] = 24'b010111110000011000111001;
rgb[14804] = 24'b011111100000100101001100;
rgb[14805] = 24'b100111100000101101011111;
rgb[14806] = 24'b101111100000110101110010;
rgb[14807] = 24'b110111100000111110000101;
rgb[14808] = 24'b111011110010000010010110;
rgb[14809] = 24'b111100010100000010100101;
rgb[14810] = 24'b111100110110000010110100;
rgb[14811] = 24'b111101011000000011000011;
rgb[14812] = 24'b111110001001111111010010;
rgb[14813] = 24'b111110101011111111100001;
rgb[14814] = 24'b111111001101111111110000;
rgb[14815] = 24'b111111111111111111111111;
rgb[14816] = 24'b000000000000000000000000;
rgb[14817] = 24'b001000000000000100010011;
rgb[14818] = 24'b010000010000001000100110;
rgb[14819] = 24'b011000100000001100111001;
rgb[14820] = 24'b100000110000010001001101;
rgb[14821] = 24'b101001000000010101100000;
rgb[14822] = 24'b110001010000011001110011;
rgb[14823] = 24'b111001100000011110000110;
rgb[14824] = 24'b111101110001100010010111;
rgb[14825] = 24'b111110000011100110100110;
rgb[14826] = 24'b111110010101101010110101;
rgb[14827] = 24'b111110100111101111000100;
rgb[14828] = 24'b111110111001110011010010;
rgb[14829] = 24'b111111001011110111100001;
rgb[14830] = 24'b111111011101111011110000;
rgb[14831] = 24'b111111111111111111111111;
rgb[14832] = 24'b000000000000000000000000;
rgb[14833] = 24'b001000100000000000010011;
rgb[14834] = 24'b010001000000000000100110;
rgb[14835] = 24'b011001100000000000111010;
rgb[14836] = 24'b100010000000000001001101;
rgb[14837] = 24'b101010100000000001100001;
rgb[14838] = 24'b110011000000000001110100;
rgb[14839] = 24'b111011100000000010001000;
rgb[14840] = 24'b111111100001000110011001;
rgb[14841] = 24'b111111110011001010100111;
rgb[14842] = 24'b111111100101010110110110;
rgb[14843] = 24'b111111110111011011000100;
rgb[14844] = 24'b111111111001100111010011;
rgb[14845] = 24'b111111111011101111100001;
rgb[14846] = 24'b111111111101110111110000;
rgb[14847] = 24'b111111111111111111111111;
rgb[14848] = 24'b000000000000000000000000;
rgb[14849] = 24'b000100010001000100010001;
rgb[14850] = 24'b001000100010001000100010;
rgb[14851] = 24'b001100110011001100110011;
rgb[14852] = 24'b010001000100010001000100;
rgb[14853] = 24'b010101010101010101010101;
rgb[14854] = 24'b011001100110011001100110;
rgb[14855] = 24'b011101110111011101110111;
rgb[14856] = 24'b100010001000100010001000;
rgb[14857] = 24'b100110011001100110011001;
rgb[14858] = 24'b101010101010101010101010;
rgb[14859] = 24'b101110111011101110111011;
rgb[14860] = 24'b110011001100110011001100;
rgb[14861] = 24'b110111011101110111011101;
rgb[14862] = 24'b111011101110111011101110;
rgb[14863] = 24'b111111111111111111111111;
rgb[14864] = 24'b000000000000000000000000;
rgb[14865] = 24'b000100100000111100010000;
rgb[14866] = 24'b001001000001111100100001;
rgb[14867] = 24'b001101100010111100110010;
rgb[14868] = 24'b010010000011111101000011;
rgb[14869] = 24'b010110100100111101010100;
rgb[14870] = 24'b011011000101111101100101;
rgb[14871] = 24'b011111100110111101110110;
rgb[14872] = 24'b100011111000000010000111;
rgb[14873] = 24'b100111111001001010011000;
rgb[14874] = 24'b101011111010010010101001;
rgb[14875] = 24'b101111111011011010111010;
rgb[14876] = 24'b110011111100100011001011;
rgb[14877] = 24'b110111111101101011011100;
rgb[14878] = 24'b111011111110110011101101;
rgb[14879] = 24'b111111111111111111111111;
rgb[14880] = 24'b000000000000000000000000;
rgb[14881] = 24'b000100110000111000010000;
rgb[14882] = 24'b001001100001110100100001;
rgb[14883] = 24'b001110010010110000110010;
rgb[14884] = 24'b010011010011101001000011;
rgb[14885] = 24'b011000000100100101010100;
rgb[14886] = 24'b011100110101100001100101;
rgb[14887] = 24'b100001100110011101110110;
rgb[14888] = 24'b100101110111100010000111;
rgb[14889] = 24'b101001101000101110011000;
rgb[14890] = 24'b101101011001111010101001;
rgb[14891] = 24'b110001001011000110111010;
rgb[14892] = 24'b110100101100010111001011;
rgb[14893] = 24'b111000011101100011011100;
rgb[14894] = 24'b111100001110101111101101;
rgb[14895] = 24'b111111111111111111111111;
rgb[14896] = 24'b000000000000000000000000;
rgb[14897] = 24'b000101000000110100010000;
rgb[14898] = 24'b001010000001101100100001;
rgb[14899] = 24'b001111010010100000110010;
rgb[14900] = 24'b010100010011011001000011;
rgb[14901] = 24'b011001010100010001010100;
rgb[14902] = 24'b011110100101000101100101;
rgb[14903] = 24'b100011100101111101110101;
rgb[14904] = 24'b100111110111000010000110;
rgb[14905] = 24'b101011011000010010011000;
rgb[14906] = 24'b101110111001100010101001;
rgb[14907] = 24'b110010001010110110111010;
rgb[14908] = 24'b110101101100000111001011;
rgb[14909] = 24'b111000111101011011011100;
rgb[14910] = 24'b111100011110101011101101;
rgb[14911] = 24'b111111111111111111111111;
rgb[14912] = 24'b000000000000000000000000;
rgb[14913] = 24'b000101010000110000010000;
rgb[14914] = 24'b001010110001100000100001;
rgb[14915] = 24'b010000000010010100110010;
rgb[14916] = 24'b010101100011000101000011;
rgb[14917] = 24'b011010110011111001010011;
rgb[14918] = 24'b100000010100101001100100;
rgb[14919] = 24'b100101100101011101110101;
rgb[14920] = 24'b101001110110100010000110;
rgb[14921] = 24'b101101000111110110010111;
rgb[14922] = 24'b110000001001001110101000;
rgb[14923] = 24'b110011011010100010111010;
rgb[14924] = 24'b110110011011111011001011;
rgb[14925] = 24'b111001101101001111011100;
rgb[14926] = 24'b111100101110100111101101;
rgb[14927] = 24'b111111111111111111111111;
rgb[14928] = 24'b000000000000000000000000;
rgb[14929] = 24'b000101100000101100010000;
rgb[14930] = 24'b001011010001011000100001;
rgb[14931] = 24'b010001000010001000110010;
rgb[14932] = 24'b010110100010110101000010;
rgb[14933] = 24'b011100010011100001010011;
rgb[14934] = 24'b100010000100010001100100;
rgb[14935] = 24'b100111100100111101110101;
rgb[14936] = 24'b101011110110000010000110;
rgb[14937] = 24'b101110110111011010010111;
rgb[14938] = 24'b110001101000110110101000;
rgb[14939] = 24'b110100011010010010111001;
rgb[14940] = 24'b110111011011101111001011;
rgb[14941] = 24'b111010001101000111011100;
rgb[14942] = 24'b111100111110100011101101;
rgb[14943] = 24'b111111111111111111111111;
rgb[14944] = 24'b000000000000000000000000;
rgb[14945] = 24'b000101110000101000010000;
rgb[14946] = 24'b001011110001010000100001;
rgb[14947] = 24'b010001110001111000110010;
rgb[14948] = 24'b010111110010100001000010;
rgb[14949] = 24'b011101100011001101010011;
rgb[14950] = 24'b100011100011110101100100;
rgb[14951] = 24'b101001100100011101110100;
rgb[14952] = 24'b101101110101100010000101;
rgb[14953] = 24'b110000010111000010010111;
rgb[14954] = 24'b110011001000011110101000;
rgb[14955] = 24'b110101101001111110111001;
rgb[14956] = 24'b111000001011011111001011;
rgb[14957] = 24'b111010101100111111011100;
rgb[14958] = 24'b111101001110011111101101;
rgb[14959] = 24'b111111101111111111111111;
rgb[14960] = 24'b000000000000000000000000;
rgb[14961] = 24'b000110000000100100010000;
rgb[14962] = 24'b001100010001001000100001;
rgb[14963] = 24'b010010100001101100110001;
rgb[14964] = 24'b011000110010010001000010;
rgb[14965] = 24'b011111000010110101010011;
rgb[14966] = 24'b100101010011011001100011;
rgb[14967] = 24'b101011100011111101110100;
rgb[14968] = 24'b101111110101000010000101;
rgb[14969] = 24'b110010000110100110010110;
rgb[14970] = 24'b110100011000001010101000;
rgb[14971] = 24'b110110101001101110111001;
rgb[14972] = 24'b111000111011010011001010;
rgb[14973] = 24'b111011001100110111011100;
rgb[14974] = 24'b111101011110011011101101;
rgb[14975] = 24'b111111111111111111111111;
rgb[14976] = 24'b000000000000000000000000;
rgb[14977] = 24'b000110100000011100010000;
rgb[14978] = 24'b001101000000111100100001;
rgb[14979] = 24'b010011100001011100110001;
rgb[14980] = 24'b011010000001111101000010;
rgb[14981] = 24'b100000100010011101010010;
rgb[14982] = 24'b100111000010111101100011;
rgb[14983] = 24'b101101100011011101110011;
rgb[14984] = 24'b110001110100100010000100;
rgb[14985] = 24'b110011110110001010010110;
rgb[14986] = 24'b110101110111110010100111;
rgb[14987] = 24'b110111111001011010111001;
rgb[14988] = 24'b111001111011000011001010;
rgb[14989] = 24'b111011111100101011011100;
rgb[14990] = 24'b111101111110010011101101;
rgb[14991] = 24'b111111101111111111111111;
rgb[14992] = 24'b000000000000000000000000;
rgb[14993] = 24'b000110110000011000010000;
rgb[14994] = 24'b001101100000110100100001;
rgb[14995] = 24'b010100010001010000110001;
rgb[14996] = 24'b011011000001101101000010;
rgb[14997] = 24'b100010000010000101010010;
rgb[14998] = 24'b101000110010100001100011;
rgb[14999] = 24'b101111100010111101110011;
rgb[15000] = 24'b110011110100000010000100;
rgb[15001] = 24'b110101100101101110010110;
rgb[15002] = 24'b110111010111011010100111;
rgb[15003] = 24'b111000111001001010111001;
rgb[15004] = 24'b111010101010110111001010;
rgb[15005] = 24'b111100011100100011011100;
rgb[15006] = 24'b111110001110001111101101;
rgb[15007] = 24'b111111111111111111111111;
rgb[15008] = 24'b000000000000000000000000;
rgb[15009] = 24'b000111000000010100010000;
rgb[15010] = 24'b001110000000101100100000;
rgb[15011] = 24'b010101010001000100110001;
rgb[15012] = 24'b011100010001011001000001;
rgb[15013] = 24'b100011010001110001010010;
rgb[15014] = 24'b101010100010001001100010;
rgb[15015] = 24'b110001100010011101110011;
rgb[15016] = 24'b110101110011100010000100;
rgb[15017] = 24'b110111010101010010010101;
rgb[15018] = 24'b111000100111000110100111;
rgb[15019] = 24'b111010001000110110111000;
rgb[15020] = 24'b111011101010101011001010;
rgb[15021] = 24'b111100111100011011011011;
rgb[15022] = 24'b111110011110001011101101;
rgb[15023] = 24'b111111101111111111111111;
rgb[15024] = 24'b000000000000000000000000;
rgb[15025] = 24'b000111010000010000010000;
rgb[15026] = 24'b001110100000100100100000;
rgb[15027] = 24'b010110000000110100110001;
rgb[15028] = 24'b011101010001001001000001;
rgb[15029] = 24'b100100110001011001010010;
rgb[15030] = 24'b101100000001101101100010;
rgb[15031] = 24'b110011100001111101110010;
rgb[15032] = 24'b110111110011000010000011;
rgb[15033] = 24'b111000110100111010010101;
rgb[15034] = 24'b111010000110101110100111;
rgb[15035] = 24'b111011001000100110111000;
rgb[15036] = 24'b111100011010011011001010;
rgb[15037] = 24'b111101011100010011011011;
rgb[15038] = 24'b111110101110000111101101;
rgb[15039] = 24'b111111111111111111111111;
rgb[15040] = 24'b000000000000000000000000;
rgb[15041] = 24'b000111100000001100010000;
rgb[15042] = 24'b001111010000011000100000;
rgb[15043] = 24'b010110110000101000110001;
rgb[15044] = 24'b011110100000110101000001;
rgb[15045] = 24'b100110010001000001010001;
rgb[15046] = 24'b101101110001010001100010;
rgb[15047] = 24'b110101100001011101110010;
rgb[15048] = 24'b111001110010100010000011;
rgb[15049] = 24'b111010100100011110010101;
rgb[15050] = 24'b111011100110010110100110;
rgb[15051] = 24'b111100011000010010111000;
rgb[15052] = 24'b111101001010001111001010;
rgb[15053] = 24'b111110001100000111011011;
rgb[15054] = 24'b111110111110000011101101;
rgb[15055] = 24'b111111111111111111111111;
rgb[15056] = 24'b000000000000000000000000;
rgb[15057] = 24'b000111110000001000010000;
rgb[15058] = 24'b001111110000010000100000;
rgb[15059] = 24'b010111110000011000110000;
rgb[15060] = 24'b011111100000100101000001;
rgb[15061] = 24'b100111100000101101010001;
rgb[15062] = 24'b101111100000110101100001;
rgb[15063] = 24'b110111100000111101110010;
rgb[15064] = 24'b111011110010000010000011;
rgb[15065] = 24'b111100010100000010010100;
rgb[15066] = 24'b111100110110000010100110;
rgb[15067] = 24'b111101011000000010111000;
rgb[15068] = 24'b111110001001111111001001;
rgb[15069] = 24'b111110101011111111011011;
rgb[15070] = 24'b111111001101111111101101;
rgb[15071] = 24'b111111111111111111111111;
rgb[15072] = 24'b000000000000000000000000;
rgb[15073] = 24'b001000000000000100010000;
rgb[15074] = 24'b010000010000001000100000;
rgb[15075] = 24'b011000100000001100110000;
rgb[15076] = 24'b100000110000010001000000;
rgb[15077] = 24'b101001000000010101010001;
rgb[15078] = 24'b110001010000011001100001;
rgb[15079] = 24'b111001100000011101110001;
rgb[15080] = 24'b111101110001100010000010;
rgb[15081] = 24'b111110000011100110010100;
rgb[15082] = 24'b111110010101101010100110;
rgb[15083] = 24'b111110100111101110110111;
rgb[15084] = 24'b111110111001110011001001;
rgb[15085] = 24'b111111001011110111011011;
rgb[15086] = 24'b111111011101111011101101;
rgb[15087] = 24'b111111111111111111111111;
rgb[15088] = 24'b000000000000000000000000;
rgb[15089] = 24'b001000100000000000010000;
rgb[15090] = 24'b010001000000000000100000;
rgb[15091] = 24'b011001100000000000110000;
rgb[15092] = 24'b100010000000000001000000;
rgb[15093] = 24'b101010100000000001010000;
rgb[15094] = 24'b110011000000000001100001;
rgb[15095] = 24'b111011100000000001110001;
rgb[15096] = 24'b111111100001000110000010;
rgb[15097] = 24'b111111110011001010010100;
rgb[15098] = 24'b111111100101010110100101;
rgb[15099] = 24'b111111110111011010110111;
rgb[15100] = 24'b111111111001100111001001;
rgb[15101] = 24'b111111111011101111011011;
rgb[15102] = 24'b111111111101110111101101;
rgb[15103] = 24'b111111111111111111111111;
rgb[15104] = 24'b000000000000000000000000;
rgb[15105] = 24'b000100010001000100010001;
rgb[15106] = 24'b001000100010001000100010;
rgb[15107] = 24'b001100110011001100110011;
rgb[15108] = 24'b010001000100010001000100;
rgb[15109] = 24'b010101010101010101010101;
rgb[15110] = 24'b011001100110011001100110;
rgb[15111] = 24'b011101110111011101110111;
rgb[15112] = 24'b100010001000100010001000;
rgb[15113] = 24'b100110011001100110011001;
rgb[15114] = 24'b101010101010101010101010;
rgb[15115] = 24'b101110111011101110111011;
rgb[15116] = 24'b110011001100110011001100;
rgb[15117] = 24'b110111011101110111011101;
rgb[15118] = 24'b111011101110111011101110;
rgb[15119] = 24'b111111111111111111111111;
rgb[15120] = 24'b000000000000000000000000;
rgb[15121] = 24'b000100100000111100010000;
rgb[15122] = 24'b001001000001111100100001;
rgb[15123] = 24'b001101100010111100110010;
rgb[15124] = 24'b010010000011111101000010;
rgb[15125] = 24'b010110100100111101010011;
rgb[15126] = 24'b011011000101111101100100;
rgb[15127] = 24'b011111100110111101110101;
rgb[15128] = 24'b100011111000000010000110;
rgb[15129] = 24'b100111111001001010010111;
rgb[15130] = 24'b101011111010010010101000;
rgb[15131] = 24'b101111111011011010111001;
rgb[15132] = 24'b110011111100100011001011;
rgb[15133] = 24'b110111111101101011011100;
rgb[15134] = 24'b111011111110110011101101;
rgb[15135] = 24'b111111111111111111111111;
rgb[15136] = 24'b000000000000000000000000;
rgb[15137] = 24'b000100110000111000010000;
rgb[15138] = 24'b001001100001110100100000;
rgb[15139] = 24'b001110010010110000110001;
rgb[15140] = 24'b010011010011101001000001;
rgb[15141] = 24'b011000000100100101010010;
rgb[15142] = 24'b011100110101100001100010;
rgb[15143] = 24'b100001100110011101110011;
rgb[15144] = 24'b100101110111100010000100;
rgb[15145] = 24'b101001101000101110010101;
rgb[15146] = 24'b101101011001111010100111;
rgb[15147] = 24'b110001001011000110111000;
rgb[15148] = 24'b110100101100010111001010;
rgb[15149] = 24'b111000011101100011011011;
rgb[15150] = 24'b111100001110101111101101;
rgb[15151] = 24'b111111111111111111111111;
rgb[15152] = 24'b000000000000000000000000;
rgb[15153] = 24'b000101000000110100010000;
rgb[15154] = 24'b001010000001101100100000;
rgb[15155] = 24'b001111010010100000110000;
rgb[15156] = 24'b010100010011011001000000;
rgb[15157] = 24'b011001010100010001010000;
rgb[15158] = 24'b011110100101000101100001;
rgb[15159] = 24'b100011100101111101110001;
rgb[15160] = 24'b100111110111000010000010;
rgb[15161] = 24'b101011011000010010010100;
rgb[15162] = 24'b101110111001100010100101;
rgb[15163] = 24'b110010001010110110110111;
rgb[15164] = 24'b110101101100000111001001;
rgb[15165] = 24'b111000111101011011011011;
rgb[15166] = 24'b111100011110101011101101;
rgb[15167] = 24'b111111111111111111111111;
rgb[15168] = 24'b000000000000000000000000;
rgb[15169] = 24'b000101010000110000001111;
rgb[15170] = 24'b001010110001100000011111;
rgb[15171] = 24'b010000000010010100101111;
rgb[15172] = 24'b010101100011000100111111;
rgb[15173] = 24'b011010110011111001001111;
rgb[15174] = 24'b100000010100101001011111;
rgb[15175] = 24'b100101100101011101101111;
rgb[15176] = 24'b101001110110100010000000;
rgb[15177] = 24'b101101000111110110010010;
rgb[15178] = 24'b110000001001001110100100;
rgb[15179] = 24'b110011011010100010110110;
rgb[15180] = 24'b110110011011111011001000;
rgb[15181] = 24'b111001101101001111011010;
rgb[15182] = 24'b111100101110100111101100;
rgb[15183] = 24'b111111111111111111111111;
rgb[15184] = 24'b000000000000000000000000;
rgb[15185] = 24'b000101100000101100001111;
rgb[15186] = 24'b001011010001011000011111;
rgb[15187] = 24'b010001000010001000101110;
rgb[15188] = 24'b010110100010110100111110;
rgb[15189] = 24'b011100010011100001001110;
rgb[15190] = 24'b100010000100010001011101;
rgb[15191] = 24'b100111100100111101101101;
rgb[15192] = 24'b101011110110000001111110;
rgb[15193] = 24'b101110110111011010010000;
rgb[15194] = 24'b110001101000110110100011;
rgb[15195] = 24'b110100011010010010110101;
rgb[15196] = 24'b110111011011101111000111;
rgb[15197] = 24'b111010001101000111011010;
rgb[15198] = 24'b111100111110100011101100;
rgb[15199] = 24'b111111111111111111111111;
rgb[15200] = 24'b000000000000000000000000;
rgb[15201] = 24'b000101110000101000001111;
rgb[15202] = 24'b001011110001010000011110;
rgb[15203] = 24'b010001110001111000101110;
rgb[15204] = 24'b010111110010100000111101;
rgb[15205] = 24'b011101100011001101001100;
rgb[15206] = 24'b100011100011110101011100;
rgb[15207] = 24'b101001100100011101101011;
rgb[15208] = 24'b101101110101100001111100;
rgb[15209] = 24'b110000010111000010001111;
rgb[15210] = 24'b110011001000011110100001;
rgb[15211] = 24'b110101101001111110110100;
rgb[15212] = 24'b111000001011011111000111;
rgb[15213] = 24'b111010101100111111011001;
rgb[15214] = 24'b111101001110011111101100;
rgb[15215] = 24'b111111101111111111111111;
rgb[15216] = 24'b000000000000000000000000;
rgb[15217] = 24'b000110000000100100001111;
rgb[15218] = 24'b001100010001001000011110;
rgb[15219] = 24'b010010100001101100101101;
rgb[15220] = 24'b011000110010010000111100;
rgb[15221] = 24'b011111000010110101001011;
rgb[15222] = 24'b100101010011011001011010;
rgb[15223] = 24'b101011100011111101101001;
rgb[15224] = 24'b101111110101000001111010;
rgb[15225] = 24'b110010000110100110001101;
rgb[15226] = 24'b110100011000001010100000;
rgb[15227] = 24'b110110101001101110110011;
rgb[15228] = 24'b111000111011010011000110;
rgb[15229] = 24'b111011001100110111011001;
rgb[15230] = 24'b111101011110011011101100;
rgb[15231] = 24'b111111111111111111111111;
rgb[15232] = 24'b000000000000000000000000;
rgb[15233] = 24'b000110100000011100001110;
rgb[15234] = 24'b001101000000111100011101;
rgb[15235] = 24'b010011100001011100101100;
rgb[15236] = 24'b011010000001111100111011;
rgb[15237] = 24'b100000100010011101001010;
rgb[15238] = 24'b100111000010111101011001;
rgb[15239] = 24'b101101100011011101100111;
rgb[15240] = 24'b110001110100100001111000;
rgb[15241] = 24'b110011110110001010001100;
rgb[15242] = 24'b110101110111110010011111;
rgb[15243] = 24'b110111111001011010110010;
rgb[15244] = 24'b111001111011000011000101;
rgb[15245] = 24'b111011111100101011011000;
rgb[15246] = 24'b111101111110010011101011;
rgb[15247] = 24'b111111101111111111111111;
rgb[15248] = 24'b000000000000000000000000;
rgb[15249] = 24'b000110110000011000001110;
rgb[15250] = 24'b001101100000110100011101;
rgb[15251] = 24'b010100010001010000101011;
rgb[15252] = 24'b011011000001101100111010;
rgb[15253] = 24'b100010000010000101001000;
rgb[15254] = 24'b101000110010100001010111;
rgb[15255] = 24'b101111100010111101100101;
rgb[15256] = 24'b110011110100000001110110;
rgb[15257] = 24'b110101100101101110001010;
rgb[15258] = 24'b110111010111011010011101;
rgb[15259] = 24'b111000111001001010110001;
rgb[15260] = 24'b111010101010110111000100;
rgb[15261] = 24'b111100011100100011011000;
rgb[15262] = 24'b111110001110001111101011;
rgb[15263] = 24'b111111111111111111111111;
rgb[15264] = 24'b000000000000000000000000;
rgb[15265] = 24'b000111000000010100001110;
rgb[15266] = 24'b001110000000101100011100;
rgb[15267] = 24'b010101010001000100101010;
rgb[15268] = 24'b011100010001011000111001;
rgb[15269] = 24'b100011010001110001000111;
rgb[15270] = 24'b101010100010001001010101;
rgb[15271] = 24'b110001100010011101100100;
rgb[15272] = 24'b110101110011100001110101;
rgb[15273] = 24'b110111010101010010001000;
rgb[15274] = 24'b111000100111000110011100;
rgb[15275] = 24'b111010001000110110110000;
rgb[15276] = 24'b111011101010101011000011;
rgb[15277] = 24'b111100111100011011010111;
rgb[15278] = 24'b111110011110001011101011;
rgb[15279] = 24'b111111101111111111111111;
rgb[15280] = 24'b000000000000000000000000;
rgb[15281] = 24'b000111010000010000001110;
rgb[15282] = 24'b001110100000100100011100;
rgb[15283] = 24'b010110000000110100101010;
rgb[15284] = 24'b011101010001001000111000;
rgb[15285] = 24'b100100110001011001000110;
rgb[15286] = 24'b101100000001101101010100;
rgb[15287] = 24'b110011100001111101100010;
rgb[15288] = 24'b110111110011000001110011;
rgb[15289] = 24'b111000110100111010000111;
rgb[15290] = 24'b111010000110101110011011;
rgb[15291] = 24'b111011001000100110101111;
rgb[15292] = 24'b111100011010011011000011;
rgb[15293] = 24'b111101011100010011010111;
rgb[15294] = 24'b111110101110000111101011;
rgb[15295] = 24'b111111111111111111111111;
rgb[15296] = 24'b000000000000000000000000;
rgb[15297] = 24'b000111100000001100001101;
rgb[15298] = 24'b001111010000011000011011;
rgb[15299] = 24'b010110110000101000101001;
rgb[15300] = 24'b011110100000110100110111;
rgb[15301] = 24'b100110010001000001000100;
rgb[15302] = 24'b101101110001010001010010;
rgb[15303] = 24'b110101100001011101100000;
rgb[15304] = 24'b111001110010100001110001;
rgb[15305] = 24'b111010100100011110000101;
rgb[15306] = 24'b111011100110010110011001;
rgb[15307] = 24'b111100011000010010101110;
rgb[15308] = 24'b111101001010001111000010;
rgb[15309] = 24'b111110001100000111010110;
rgb[15310] = 24'b111110111110000011101010;
rgb[15311] = 24'b111111111111111111111111;
rgb[15312] = 24'b000000000000000000000000;
rgb[15313] = 24'b000111110000001000001101;
rgb[15314] = 24'b001111110000010000011010;
rgb[15315] = 24'b010111110000011000101000;
rgb[15316] = 24'b011111100000100100110101;
rgb[15317] = 24'b100111100000101101000011;
rgb[15318] = 24'b101111100000110101010000;
rgb[15319] = 24'b110111100000111101011110;
rgb[15320] = 24'b111011110010000001101111;
rgb[15321] = 24'b111100010100000010000011;
rgb[15322] = 24'b111100110110000010011000;
rgb[15323] = 24'b111101011000000010101100;
rgb[15324] = 24'b111110001001111111000001;
rgb[15325] = 24'b111110101011111111010101;
rgb[15326] = 24'b111111001101111111101010;
rgb[15327] = 24'b111111111111111111111111;
rgb[15328] = 24'b000000000000000000000000;
rgb[15329] = 24'b001000000000000100001101;
rgb[15330] = 24'b010000010000001000011010;
rgb[15331] = 24'b011000100000001100100111;
rgb[15332] = 24'b100000110000010000110100;
rgb[15333] = 24'b101001000000010101000010;
rgb[15334] = 24'b110001010000011001001111;
rgb[15335] = 24'b111001100000011101011100;
rgb[15336] = 24'b111101110001100001101101;
rgb[15337] = 24'b111110000011100110000010;
rgb[15338] = 24'b111110010101101010010111;
rgb[15339] = 24'b111110100111101110101011;
rgb[15340] = 24'b111110111001110011000000;
rgb[15341] = 24'b111111001011110111010101;
rgb[15342] = 24'b111111011101111011101010;
rgb[15343] = 24'b111111111111111111111111;
rgb[15344] = 24'b000000000000000000000000;
rgb[15345] = 24'b001000100000000000001100;
rgb[15346] = 24'b010001000000000000011001;
rgb[15347] = 24'b011001100000000000100110;
rgb[15348] = 24'b100010000000000000110011;
rgb[15349] = 24'b101010100000000001000000;
rgb[15350] = 24'b110011000000000001001101;
rgb[15351] = 24'b111011100000000001011010;
rgb[15352] = 24'b111111100001000101101011;
rgb[15353] = 24'b111111110011001010000000;
rgb[15354] = 24'b111111100101010110010101;
rgb[15355] = 24'b111111110111011010101010;
rgb[15356] = 24'b111111111001100110111111;
rgb[15357] = 24'b111111111011101111010100;
rgb[15358] = 24'b111111111101110111101001;
rgb[15359] = 24'b111111111111111111111111;
rgb[15360] = 24'b000000000000000000000000;
rgb[15361] = 24'b000100010001000100010001;
rgb[15362] = 24'b001000100010001000100010;
rgb[15363] = 24'b001100110011001100110011;
rgb[15364] = 24'b010001000100010001000100;
rgb[15365] = 24'b010101010101010101010101;
rgb[15366] = 24'b011001100110011001100110;
rgb[15367] = 24'b011101110111011101110111;
rgb[15368] = 24'b100010001000100010001000;
rgb[15369] = 24'b100110011001100110011001;
rgb[15370] = 24'b101010101010101010101010;
rgb[15371] = 24'b101110111011101110111011;
rgb[15372] = 24'b110011001100110011001100;
rgb[15373] = 24'b110111011101110111011101;
rgb[15374] = 24'b111011101110111011101110;
rgb[15375] = 24'b111111111111111111111111;
rgb[15376] = 24'b000000000000000000000000;
rgb[15377] = 24'b000100100000111100010000;
rgb[15378] = 24'b001001000001111100100001;
rgb[15379] = 24'b001101100010111100110001;
rgb[15380] = 24'b010010000011111101000010;
rgb[15381] = 24'b010110100100111101010010;
rgb[15382] = 24'b011011000101111101100011;
rgb[15383] = 24'b011111100110111101110011;
rgb[15384] = 24'b100011111000000010000100;
rgb[15385] = 24'b100111111001001010010110;
rgb[15386] = 24'b101011111010010010100111;
rgb[15387] = 24'b101111111011011010111001;
rgb[15388] = 24'b110011111100100011001010;
rgb[15389] = 24'b110111111101101011011100;
rgb[15390] = 24'b111011111110110011101101;
rgb[15391] = 24'b111111111111111111111111;
rgb[15392] = 24'b000000000000000000000000;
rgb[15393] = 24'b000100110000111000010000;
rgb[15394] = 24'b001001100001110100100000;
rgb[15395] = 24'b001110010010110000110000;
rgb[15396] = 24'b010011010011101001000000;
rgb[15397] = 24'b011000000100100101010000;
rgb[15398] = 24'b011100110101100001100000;
rgb[15399] = 24'b100001100110011101110000;
rgb[15400] = 24'b100101110111100010000001;
rgb[15401] = 24'b101001101000101110010011;
rgb[15402] = 24'b101101011001111010100101;
rgb[15403] = 24'b110001001011000110110111;
rgb[15404] = 24'b110100101100010111001001;
rgb[15405] = 24'b111000011101100011011011;
rgb[15406] = 24'b111100001110101111101101;
rgb[15407] = 24'b111111111111111111111111;
rgb[15408] = 24'b000000000000000000000000;
rgb[15409] = 24'b000101000000110100001111;
rgb[15410] = 24'b001010000001101100011111;
rgb[15411] = 24'b001111010010100000101110;
rgb[15412] = 24'b010100010011011000111110;
rgb[15413] = 24'b011001010100010001001101;
rgb[15414] = 24'b011110100101000101011101;
rgb[15415] = 24'b100011100101111101101100;
rgb[15416] = 24'b100111110111000001111101;
rgb[15417] = 24'b101011011000010010010000;
rgb[15418] = 24'b101110111001100010100010;
rgb[15419] = 24'b110010001010110110110101;
rgb[15420] = 24'b110101101100000111000111;
rgb[15421] = 24'b111000111101011011011010;
rgb[15422] = 24'b111100011110101011101100;
rgb[15423] = 24'b111111111111111111111111;
rgb[15424] = 24'b000000000000000000000000;
rgb[15425] = 24'b000101010000110000001111;
rgb[15426] = 24'b001010110001100000011110;
rgb[15427] = 24'b010000000010010100101101;
rgb[15428] = 24'b010101100011000100111100;
rgb[15429] = 24'b011010110011111001001011;
rgb[15430] = 24'b100000010100101001011010;
rgb[15431] = 24'b100101100101011101101001;
rgb[15432] = 24'b101001110110100001111010;
rgb[15433] = 24'b101101000111110110001101;
rgb[15434] = 24'b110000001001001110100000;
rgb[15435] = 24'b110011011010100010110011;
rgb[15436] = 24'b110110011011111011000110;
rgb[15437] = 24'b111001101101001111011001;
rgb[15438] = 24'b111100101110100111101100;
rgb[15439] = 24'b111111111111111111111111;
rgb[15440] = 24'b000000000000000000000000;
rgb[15441] = 24'b000101100000101100001110;
rgb[15442] = 24'b001011010001011000011101;
rgb[15443] = 24'b010001000010001000101011;
rgb[15444] = 24'b010110100010110100111010;
rgb[15445] = 24'b011100010011100001001000;
rgb[15446] = 24'b100010000100010001010111;
rgb[15447] = 24'b100111100100111101100101;
rgb[15448] = 24'b101011110110000001110110;
rgb[15449] = 24'b101110110111011010001010;
rgb[15450] = 24'b110001101000110110011101;
rgb[15451] = 24'b110100011010010010110001;
rgb[15452] = 24'b110111011011101111000100;
rgb[15453] = 24'b111010001101000111011000;
rgb[15454] = 24'b111100111110100011101011;
rgb[15455] = 24'b111111111111111111111111;
rgb[15456] = 24'b000000000000000000000000;
rgb[15457] = 24'b000101110000101000001110;
rgb[15458] = 24'b001011110001010000011100;
rgb[15459] = 24'b010001110001111000101010;
rgb[15460] = 24'b010111110010100000111000;
rgb[15461] = 24'b011101100011001101000110;
rgb[15462] = 24'b100011100011110101010100;
rgb[15463] = 24'b101001100100011101100010;
rgb[15464] = 24'b101101110101100001110011;
rgb[15465] = 24'b110000010111000010000111;
rgb[15466] = 24'b110011001000011110011011;
rgb[15467] = 24'b110101101001111110101111;
rgb[15468] = 24'b111000001011011111000011;
rgb[15469] = 24'b111010101100111111010111;
rgb[15470] = 24'b111101001110011111101011;
rgb[15471] = 24'b111111101111111111111111;
rgb[15472] = 24'b000000000000000000000000;
rgb[15473] = 24'b000110000000100100001101;
rgb[15474] = 24'b001100010001001000011011;
rgb[15475] = 24'b010010100001101100101000;
rgb[15476] = 24'b011000110010010000110110;
rgb[15477] = 24'b011111000010110101000011;
rgb[15478] = 24'b100101010011011001010001;
rgb[15479] = 24'b101011100011111101011111;
rgb[15480] = 24'b101111110101000001110000;
rgb[15481] = 24'b110010000110100110000100;
rgb[15482] = 24'b110100011000001010011000;
rgb[15483] = 24'b110110101001101110101101;
rgb[15484] = 24'b111000111011010011000001;
rgb[15485] = 24'b111011001100110111010110;
rgb[15486] = 24'b111101011110011011101010;
rgb[15487] = 24'b111111111111111111111111;
rgb[15488] = 24'b000000000000000000000000;
rgb[15489] = 24'b000110100000011100001101;
rgb[15490] = 24'b001101000000111100011010;
rgb[15491] = 24'b010011100001011100100111;
rgb[15492] = 24'b011010000001111100110100;
rgb[15493] = 24'b100000100010011101000001;
rgb[15494] = 24'b100111000010111101001110;
rgb[15495] = 24'b101101100011011101011011;
rgb[15496] = 24'b110001110100100001101100;
rgb[15497] = 24'b110011110110001010000001;
rgb[15498] = 24'b110101110111110010010110;
rgb[15499] = 24'b110111111001011010101011;
rgb[15500] = 24'b111001111011000011000000;
rgb[15501] = 24'b111011111100101011010101;
rgb[15502] = 24'b111101111110010011101010;
rgb[15503] = 24'b111111101111111111111111;
rgb[15504] = 24'b000000000000000000000000;
rgb[15505] = 24'b000110110000011000001100;
rgb[15506] = 24'b001101100000110100011001;
rgb[15507] = 24'b010100010001010000100101;
rgb[15508] = 24'b011011000001101100110010;
rgb[15509] = 24'b100010000010000100111111;
rgb[15510] = 24'b101000110010100001001011;
rgb[15511] = 24'b101111100010111101011000;
rgb[15512] = 24'b110011110100000001101001;
rgb[15513] = 24'b110101100101101101111110;
rgb[15514] = 24'b110111010111011010010100;
rgb[15515] = 24'b111000111001001010101001;
rgb[15516] = 24'b111010101010110110111110;
rgb[15517] = 24'b111100011100100011010100;
rgb[15518] = 24'b111110001110001111101001;
rgb[15519] = 24'b111111111111111111111111;
rgb[15520] = 24'b000000000000000000000000;
rgb[15521] = 24'b000111000000010100001100;
rgb[15522] = 24'b001110000000101100011000;
rgb[15523] = 24'b010101010001000100100100;
rgb[15524] = 24'b011100010001011000110000;
rgb[15525] = 24'b100011010001110000111100;
rgb[15526] = 24'b101010100010001001001000;
rgb[15527] = 24'b110001100010011101010100;
rgb[15528] = 24'b110101110011100001100101;
rgb[15529] = 24'b110111010101010001111011;
rgb[15530] = 24'b111000100111000110010001;
rgb[15531] = 24'b111010001000110110100111;
rgb[15532] = 24'b111011101010101010111101;
rgb[15533] = 24'b111100111100011011010011;
rgb[15534] = 24'b111110011110001011101001;
rgb[15535] = 24'b111111101111111111111111;
rgb[15536] = 24'b000000000000000000000000;
rgb[15537] = 24'b000111010000010000001011;
rgb[15538] = 24'b001110100000100100010111;
rgb[15539] = 24'b010110000000110100100010;
rgb[15540] = 24'b011101010001001000101110;
rgb[15541] = 24'b100100110001011000111010;
rgb[15542] = 24'b101100000001101101000101;
rgb[15543] = 24'b110011100001111101010001;
rgb[15544] = 24'b110111110011000001100010;
rgb[15545] = 24'b111000110100111001111000;
rgb[15546] = 24'b111010000110101110001111;
rgb[15547] = 24'b111011001000100110100101;
rgb[15548] = 24'b111100011010011010111011;
rgb[15549] = 24'b111101011100010011010010;
rgb[15550] = 24'b111110101110000111101000;
rgb[15551] = 24'b111111111111111111111111;
rgb[15552] = 24'b000000000000000000000000;
rgb[15553] = 24'b000111100000001100001011;
rgb[15554] = 24'b001111010000011000010110;
rgb[15555] = 24'b010110110000101000100001;
rgb[15556] = 24'b011110100000110100101100;
rgb[15557] = 24'b100110010001000000110111;
rgb[15558] = 24'b101101110001010001000011;
rgb[15559] = 24'b110101100001011101001110;
rgb[15560] = 24'b111001110010100001011111;
rgb[15561] = 24'b111010100100011101110110;
rgb[15562] = 24'b111011100110010110001100;
rgb[15563] = 24'b111100011000010010100011;
rgb[15564] = 24'b111101001010001110111010;
rgb[15565] = 24'b111110001100000111010001;
rgb[15566] = 24'b111110111110000011101000;
rgb[15567] = 24'b111111111111111111111111;
rgb[15568] = 24'b000000000000000000000000;
rgb[15569] = 24'b000111110000001000001010;
rgb[15570] = 24'b001111110000010000010101;
rgb[15571] = 24'b010111110000011000100000;
rgb[15572] = 24'b011111100000100100101010;
rgb[15573] = 24'b100111100000101100110101;
rgb[15574] = 24'b101111100000110101000000;
rgb[15575] = 24'b110111100000111101001010;
rgb[15576] = 24'b111011110010000001011011;
rgb[15577] = 24'b111100010100000001110011;
rgb[15578] = 24'b111100110110000010001010;
rgb[15579] = 24'b111101011000000010100001;
rgb[15580] = 24'b111110001001111110111001;
rgb[15581] = 24'b111110101011111111010000;
rgb[15582] = 24'b111111001101111111100111;
rgb[15583] = 24'b111111111111111111111111;
rgb[15584] = 24'b000000000000000000000000;
rgb[15585] = 24'b001000000000000100001010;
rgb[15586] = 24'b010000010000001000010100;
rgb[15587] = 24'b011000100000001100011110;
rgb[15588] = 24'b100000110000010000101000;
rgb[15589] = 24'b101001000000010100110010;
rgb[15590] = 24'b110001010000011000111101;
rgb[15591] = 24'b111001100000011101000111;
rgb[15592] = 24'b111101110001100001011000;
rgb[15593] = 24'b111110000011100101110000;
rgb[15594] = 24'b111110010101101010000111;
rgb[15595] = 24'b111110100111101110011111;
rgb[15596] = 24'b111110111001110010110111;
rgb[15597] = 24'b111111001011110111001111;
rgb[15598] = 24'b111111011101111011100111;
rgb[15599] = 24'b111111111111111111111111;
rgb[15600] = 24'b000000000000000000000000;
rgb[15601] = 24'b001000100000000000001001;
rgb[15602] = 24'b010001000000000000010011;
rgb[15603] = 24'b011001100000000000011101;
rgb[15604] = 24'b100010000000000000100110;
rgb[15605] = 24'b101010100000000000110000;
rgb[15606] = 24'b110011000000000000111010;
rgb[15607] = 24'b111011100000000001000011;
rgb[15608] = 24'b111111100001000101010100;
rgb[15609] = 24'b111111110011001001101101;
rgb[15610] = 24'b111111100101010110000101;
rgb[15611] = 24'b111111110111011010011101;
rgb[15612] = 24'b111111111001100110110110;
rgb[15613] = 24'b111111111011101111001110;
rgb[15614] = 24'b111111111101110111100110;
rgb[15615] = 24'b111111111111111111111111;
rgb[15616] = 24'b000000000000000000000000;
rgb[15617] = 24'b000100010001000100010001;
rgb[15618] = 24'b001000100010001000100010;
rgb[15619] = 24'b001100110011001100110011;
rgb[15620] = 24'b010001000100010001000100;
rgb[15621] = 24'b010101010101010101010101;
rgb[15622] = 24'b011001100110011001100110;
rgb[15623] = 24'b011101110111011101110111;
rgb[15624] = 24'b100010001000100010001000;
rgb[15625] = 24'b100110011001100110011001;
rgb[15626] = 24'b101010101010101010101010;
rgb[15627] = 24'b101110111011101110111011;
rgb[15628] = 24'b110011001100110011001100;
rgb[15629] = 24'b110111011101110111011101;
rgb[15630] = 24'b111011101110111011101110;
rgb[15631] = 24'b111111111111111111111111;
rgb[15632] = 24'b000000000000000000000000;
rgb[15633] = 24'b000100100000111100010000;
rgb[15634] = 24'b001001000001111100100000;
rgb[15635] = 24'b001101100010111100110000;
rgb[15636] = 24'b010010000011111101000001;
rgb[15637] = 24'b010110100100111101010001;
rgb[15638] = 24'b011011000101111101100001;
rgb[15639] = 24'b011111100110111101110010;
rgb[15640] = 24'b100011111000000010000011;
rgb[15641] = 24'b100111111001001010010100;
rgb[15642] = 24'b101011111010010010100110;
rgb[15643] = 24'b101111111011011010111000;
rgb[15644] = 24'b110011111100100011001001;
rgb[15645] = 24'b110111111101101011011011;
rgb[15646] = 24'b111011111110110011101101;
rgb[15647] = 24'b111111111111111111111111;
rgb[15648] = 24'b000000000000000000000000;
rgb[15649] = 24'b000100110000111000001111;
rgb[15650] = 24'b001001100001110100011111;
rgb[15651] = 24'b001110010010110000101110;
rgb[15652] = 24'b010011010011101000111110;
rgb[15653] = 24'b011000000100100101001101;
rgb[15654] = 24'b011100110101100001011101;
rgb[15655] = 24'b100001100110011101101101;
rgb[15656] = 24'b100101110111100001111110;
rgb[15657] = 24'b101001101000101110010000;
rgb[15658] = 24'b101101011001111010100010;
rgb[15659] = 24'b110001001011000110110101;
rgb[15660] = 24'b110100101100010111000111;
rgb[15661] = 24'b111000011101100011011010;
rgb[15662] = 24'b111100001110101111101100;
rgb[15663] = 24'b111111111111111111111111;
rgb[15664] = 24'b000000000000000000000000;
rgb[15665] = 24'b000101000000110100001110;
rgb[15666] = 24'b001010000001101100011101;
rgb[15667] = 24'b001111010010100000101100;
rgb[15668] = 24'b010100010011011000111011;
rgb[15669] = 24'b011001010100010001001010;
rgb[15670] = 24'b011110100101000101011001;
rgb[15671] = 24'b100011100101111101101000;
rgb[15672] = 24'b100111110111000001111001;
rgb[15673] = 24'b101011011000010010001100;
rgb[15674] = 24'b101110111001100010011111;
rgb[15675] = 24'b110010001010110110110010;
rgb[15676] = 24'b110101101100000111000101;
rgb[15677] = 24'b111000111101011011011000;
rgb[15678] = 24'b111100011110101011101011;
rgb[15679] = 24'b111111111111111111111111;
rgb[15680] = 24'b000000000000000000000000;
rgb[15681] = 24'b000101010000110000001110;
rgb[15682] = 24'b001010110001100000011100;
rgb[15683] = 24'b010000000010010100101010;
rgb[15684] = 24'b010101100011000100111000;
rgb[15685] = 24'b011010110011111001000110;
rgb[15686] = 24'b100000010100101001010101;
rgb[15687] = 24'b100101100101011101100011;
rgb[15688] = 24'b101001110110100001110100;
rgb[15689] = 24'b101101000111110110001000;
rgb[15690] = 24'b110000001001001110011011;
rgb[15691] = 24'b110011011010100010101111;
rgb[15692] = 24'b110110011011111011000011;
rgb[15693] = 24'b111001101101001111010111;
rgb[15694] = 24'b111100101110100111101011;
rgb[15695] = 24'b111111111111111111111111;
rgb[15696] = 24'b000000000000000000000000;
rgb[15697] = 24'b000101100000101100001101;
rgb[15698] = 24'b001011010001011000011010;
rgb[15699] = 24'b010001000010001000101000;
rgb[15700] = 24'b010110100010110100110101;
rgb[15701] = 24'b011100010011100001000011;
rgb[15702] = 24'b100010000100010001010000;
rgb[15703] = 24'b100111100100111101011110;
rgb[15704] = 24'b101011110110000001101111;
rgb[15705] = 24'b101110110111011010000011;
rgb[15706] = 24'b110001101000110110011000;
rgb[15707] = 24'b110100011010010010101100;
rgb[15708] = 24'b110111011011101111000001;
rgb[15709] = 24'b111010001101000111010101;
rgb[15710] = 24'b111100111110100011101010;
rgb[15711] = 24'b111111111111111111111111;
rgb[15712] = 24'b000000000000000000000000;
rgb[15713] = 24'b000101110000101000001100;
rgb[15714] = 24'b001011110001010000011001;
rgb[15715] = 24'b010001110001111000100110;
rgb[15716] = 24'b010111110010100000110011;
rgb[15717] = 24'b011101100011001100111111;
rgb[15718] = 24'b100011100011110101001100;
rgb[15719] = 24'b101001100100011101011001;
rgb[15720] = 24'b101101110101100001101010;
rgb[15721] = 24'b110000010111000001111111;
rgb[15722] = 24'b110011001000011110010100;
rgb[15723] = 24'b110101101001111110101010;
rgb[15724] = 24'b111000001011011110111111;
rgb[15725] = 24'b111010101100111111010100;
rgb[15726] = 24'b111101001110011111101001;
rgb[15727] = 24'b111111101111111111111111;
rgb[15728] = 24'b000000000000000000000000;
rgb[15729] = 24'b000110000000100100001100;
rgb[15730] = 24'b001100010001001000011000;
rgb[15731] = 24'b010010100001101100100100;
rgb[15732] = 24'b011000110010010000110000;
rgb[15733] = 24'b011111000010110100111100;
rgb[15734] = 24'b100101010011011001001000;
rgb[15735] = 24'b101011100011111101010100;
rgb[15736] = 24'b101111110101000001100101;
rgb[15737] = 24'b110010000110100101111011;
rgb[15738] = 24'b110100011000001010010001;
rgb[15739] = 24'b110110101001101110100111;
rgb[15740] = 24'b111000111011010010111101;
rgb[15741] = 24'b111011001100110111010011;
rgb[15742] = 24'b111101011110011011101001;
rgb[15743] = 24'b111111111111111111111111;
rgb[15744] = 24'b000000000000000000000000;
rgb[15745] = 24'b000110100000011100001011;
rgb[15746] = 24'b001101000000111100010110;
rgb[15747] = 24'b010011100001011100100010;
rgb[15748] = 24'b011010000001111100101101;
rgb[15749] = 24'b100000100010011100111000;
rgb[15750] = 24'b100111000010111101000100;
rgb[15751] = 24'b101101100011011101001111;
rgb[15752] = 24'b110001110100100001100000;
rgb[15753] = 24'b110011110110001001110111;
rgb[15754] = 24'b110101110111110010001101;
rgb[15755] = 24'b110111111001011010100100;
rgb[15756] = 24'b111001111011000010111011;
rgb[15757] = 24'b111011111100101011010001;
rgb[15758] = 24'b111101111110010011101000;
rgb[15759] = 24'b111111101111111111111111;
rgb[15760] = 24'b000000000000000000000000;
rgb[15761] = 24'b000110110000011000001010;
rgb[15762] = 24'b001101100000110100010101;
rgb[15763] = 24'b010100010001010000100000;
rgb[15764] = 24'b011011000001101100101010;
rgb[15765] = 24'b100010000010000100110101;
rgb[15766] = 24'b101000110010100001000000;
rgb[15767] = 24'b101111100010111101001010;
rgb[15768] = 24'b110011110100000001011011;
rgb[15769] = 24'b110101100101101101110011;
rgb[15770] = 24'b110111010111011010001010;
rgb[15771] = 24'b111000111001001010100001;
rgb[15772] = 24'b111010101010110110111001;
rgb[15773] = 24'b111100011100100011010000;
rgb[15774] = 24'b111110001110001111100111;
rgb[15775] = 24'b111111111111111111111111;
rgb[15776] = 24'b000000000000000000000000;
rgb[15777] = 24'b000111000000010100001001;
rgb[15778] = 24'b001110000000101100010011;
rgb[15779] = 24'b010101010001000100011101;
rgb[15780] = 24'b011100010001011000100111;
rgb[15781] = 24'b100011010001110000110001;
rgb[15782] = 24'b101010100010001000111011;
rgb[15783] = 24'b110001100010011101000101;
rgb[15784] = 24'b110101110011100001010110;
rgb[15785] = 24'b110111010101010001101110;
rgb[15786] = 24'b111000100111000110000110;
rgb[15787] = 24'b111010001000110110011110;
rgb[15788] = 24'b111011101010101010110110;
rgb[15789] = 24'b111100111100011011001110;
rgb[15790] = 24'b111110011110001011100110;
rgb[15791] = 24'b111111101111111111111111;
rgb[15792] = 24'b000000000000000000000000;
rgb[15793] = 24'b000111010000010000001001;
rgb[15794] = 24'b001110100000100100010010;
rgb[15795] = 24'b010110000000110100011011;
rgb[15796] = 24'b011101010001001000100101;
rgb[15797] = 24'b100100110001011000101110;
rgb[15798] = 24'b101100000001101100110111;
rgb[15799] = 24'b110011100001111101000000;
rgb[15800] = 24'b110111110011000001010001;
rgb[15801] = 24'b111000110100111001101010;
rgb[15802] = 24'b111010000110101110000011;
rgb[15803] = 24'b111011001000100110011100;
rgb[15804] = 24'b111100011010011010110100;
rgb[15805] = 24'b111101011100010011001101;
rgb[15806] = 24'b111110101110000111100110;
rgb[15807] = 24'b111111111111111111111111;
rgb[15808] = 24'b000000000000000000000000;
rgb[15809] = 24'b000111100000001100001000;
rgb[15810] = 24'b001111010000011000010001;
rgb[15811] = 24'b010110110000101000011001;
rgb[15812] = 24'b011110100000110100100010;
rgb[15813] = 24'b100110010001000000101010;
rgb[15814] = 24'b101101110001010000110011;
rgb[15815] = 24'b110101100001011100111100;
rgb[15816] = 24'b111001110010100001001101;
rgb[15817] = 24'b111010100100011101100110;
rgb[15818] = 24'b111011100110010101111111;
rgb[15819] = 24'b111100011000010010011001;
rgb[15820] = 24'b111101001010001110110010;
rgb[15821] = 24'b111110001100000111001100;
rgb[15822] = 24'b111110111110000011100101;
rgb[15823] = 24'b111111111111111111111111;
rgb[15824] = 24'b000000000000000000000000;
rgb[15825] = 24'b000111110000001000000111;
rgb[15826] = 24'b001111110000010000001111;
rgb[15827] = 24'b010111110000011000010111;
rgb[15828] = 24'b011111100000100100011111;
rgb[15829] = 24'b100111100000101100100111;
rgb[15830] = 24'b101111100000110100101111;
rgb[15831] = 24'b110111100000111100110111;
rgb[15832] = 24'b111011110010000001001000;
rgb[15833] = 24'b111100010100000001100010;
rgb[15834] = 24'b111100110110000001111100;
rgb[15835] = 24'b111101011000000010010110;
rgb[15836] = 24'b111110001001111110110000;
rgb[15837] = 24'b111110101011111111001010;
rgb[15838] = 24'b111111001101111111100100;
rgb[15839] = 24'b111111111111111111111111;
rgb[15840] = 24'b000000000000000000000000;
rgb[15841] = 24'b001000000000000100000111;
rgb[15842] = 24'b010000010000001000001110;
rgb[15843] = 24'b011000100000001100010101;
rgb[15844] = 24'b100000110000010000011100;
rgb[15845] = 24'b101001000000010100100011;
rgb[15846] = 24'b110001010000011000101011;
rgb[15847] = 24'b111001100000011100110010;
rgb[15848] = 24'b111101110001100001000011;
rgb[15849] = 24'b111110000011100101011110;
rgb[15850] = 24'b111110010101101001111000;
rgb[15851] = 24'b111110100111101110010011;
rgb[15852] = 24'b111110111001110010101110;
rgb[15853] = 24'b111111001011110111001001;
rgb[15854] = 24'b111111011101111011100100;
rgb[15855] = 24'b111111111111111111111111;
rgb[15856] = 24'b000000000000000000000000;
rgb[15857] = 24'b001000100000000000000110;
rgb[15858] = 24'b010001000000000000001100;
rgb[15859] = 24'b011001100000000000010011;
rgb[15860] = 24'b100010000000000000011001;
rgb[15861] = 24'b101010100000000000100000;
rgb[15862] = 24'b110011000000000000100110;
rgb[15863] = 24'b111011100000000000101101;
rgb[15864] = 24'b111111100001000100111110;
rgb[15865] = 24'b111111110011001001011001;
rgb[15866] = 24'b111111100101010101110101;
rgb[15867] = 24'b111111110111011010010000;
rgb[15868] = 24'b111111111001100110101100;
rgb[15869] = 24'b111111111011101111000111;
rgb[15870] = 24'b111111111101110111100011;
rgb[15871] = 24'b111111111111111111111111;
rgb[15872] = 24'b000000000000000000000000;
rgb[15873] = 24'b000100010001000100010001;
rgb[15874] = 24'b001000100010001000100010;
rgb[15875] = 24'b001100110011001100110011;
rgb[15876] = 24'b010001000100010001000100;
rgb[15877] = 24'b010101010101010101010101;
rgb[15878] = 24'b011001100110011001100110;
rgb[15879] = 24'b011101110111011101110111;
rgb[15880] = 24'b100010001000100010001000;
rgb[15881] = 24'b100110011001100110011001;
rgb[15882] = 24'b101010101010101010101010;
rgb[15883] = 24'b101110111011101110111011;
rgb[15884] = 24'b110011001100110011001100;
rgb[15885] = 24'b110111011101110111011101;
rgb[15886] = 24'b111011101110111011101110;
rgb[15887] = 24'b111111111111111111111111;
rgb[15888] = 24'b000000000000000000000000;
rgb[15889] = 24'b000100100000111100010000;
rgb[15890] = 24'b001001000001111100100000;
rgb[15891] = 24'b001101100010111100110000;
rgb[15892] = 24'b010010000011111101000000;
rgb[15893] = 24'b010110100100111101010000;
rgb[15894] = 24'b011011000101111101100000;
rgb[15895] = 24'b011111100110111101110000;
rgb[15896] = 24'b100011111000000010000001;
rgb[15897] = 24'b100111111001001010010011;
rgb[15898] = 24'b101011111010010010100101;
rgb[15899] = 24'b101111111011011010110111;
rgb[15900] = 24'b110011111100100011001001;
rgb[15901] = 24'b110111111101101011011011;
rgb[15902] = 24'b111011111110110011101101;
rgb[15903] = 24'b111111111111111111111111;
rgb[15904] = 24'b000000000000000000000000;
rgb[15905] = 24'b000100110000111000001111;
rgb[15906] = 24'b001001100001110100011110;
rgb[15907] = 24'b001110010010110000101101;
rgb[15908] = 24'b010011010011101000111100;
rgb[15909] = 24'b011000000100100101001011;
rgb[15910] = 24'b011100110101100001011010;
rgb[15911] = 24'b100001100110011101101010;
rgb[15912] = 24'b100101110111100001111011;
rgb[15913] = 24'b101001101000101110001101;
rgb[15914] = 24'b101101011001111010100000;
rgb[15915] = 24'b110001001011000110110011;
rgb[15916] = 24'b110100101100010111000110;
rgb[15917] = 24'b111000011101100011011001;
rgb[15918] = 24'b111100001110101111101100;
rgb[15919] = 24'b111111111111111111111111;
rgb[15920] = 24'b000000000000000000000000;
rgb[15921] = 24'b000101000000110100001110;
rgb[15922] = 24'b001010000001101100011100;
rgb[15923] = 24'b001111010010100000101010;
rgb[15924] = 24'b010100010011011000111000;
rgb[15925] = 24'b011001010100010001000111;
rgb[15926] = 24'b011110100101000101010101;
rgb[15927] = 24'b100011100101111101100011;
rgb[15928] = 24'b100111110111000001110100;
rgb[15929] = 24'b101011011000010010001000;
rgb[15930] = 24'b101110111001100010011100;
rgb[15931] = 24'b110010001010110110101111;
rgb[15932] = 24'b110101101100000111000011;
rgb[15933] = 24'b111000111101011011010111;
rgb[15934] = 24'b111100011110101011101011;
rgb[15935] = 24'b111111111111111111111111;
rgb[15936] = 24'b000000000000000000000000;
rgb[15937] = 24'b000101010000110000001101;
rgb[15938] = 24'b001010110001100000011010;
rgb[15939] = 24'b010000000010010100100111;
rgb[15940] = 24'b010101100011000100110101;
rgb[15941] = 24'b011010110011111001000010;
rgb[15942] = 24'b100000010100101001001111;
rgb[15943] = 24'b100101100101011101011101;
rgb[15944] = 24'b101001110110100001101110;
rgb[15945] = 24'b101101000111110110000010;
rgb[15946] = 24'b110000001001001110010111;
rgb[15947] = 24'b110011011010100010101100;
rgb[15948] = 24'b110110011011111011000000;
rgb[15949] = 24'b111001101101001111010101;
rgb[15950] = 24'b111100101110100111101010;
rgb[15951] = 24'b111111111111111111111111;
rgb[15952] = 24'b000000000000000000000000;
rgb[15953] = 24'b000101100000101100001100;
rgb[15954] = 24'b001011010001011000011000;
rgb[15955] = 24'b010001000010001000100101;
rgb[15956] = 24'b010110100010110100110001;
rgb[15957] = 24'b011100010011100000111110;
rgb[15958] = 24'b100010000100010001001010;
rgb[15959] = 24'b100111100100111101010110;
rgb[15960] = 24'b101011110110000001100111;
rgb[15961] = 24'b101110110111011001111101;
rgb[15962] = 24'b110001101000110110010011;
rgb[15963] = 24'b110100011010010010101000;
rgb[15964] = 24'b110111011011101110111110;
rgb[15965] = 24'b111010001101000111010011;
rgb[15966] = 24'b111100111110100011101001;
rgb[15967] = 24'b111111111111111111111111;
rgb[15968] = 24'b000000000000000000000000;
rgb[15969] = 24'b000101110000101000001011;
rgb[15970] = 24'b001011110001010000010110;
rgb[15971] = 24'b010001110001111000100010;
rgb[15972] = 24'b010111110010100000101101;
rgb[15973] = 24'b011101100011001100111001;
rgb[15974] = 24'b100011100011110101000100;
rgb[15975] = 24'b101001100100011101010000;
rgb[15976] = 24'b101101110101100001100001;
rgb[15977] = 24'b110000010111000001110111;
rgb[15978] = 24'b110011001000011110001110;
rgb[15979] = 24'b110101101001111110100100;
rgb[15980] = 24'b111000001011011110111011;
rgb[15981] = 24'b111010101100111111010001;
rgb[15982] = 24'b111101001110011111101000;
rgb[15983] = 24'b111111101111111111111111;
rgb[15984] = 24'b000000000000000000000000;
rgb[15985] = 24'b000110000000100100001010;
rgb[15986] = 24'b001100010001001000010101;
rgb[15987] = 24'b010010100001101100011111;
rgb[15988] = 24'b011000110010010000101010;
rgb[15989] = 24'b011111000010110100110100;
rgb[15990] = 24'b100101010011011000111111;
rgb[15991] = 24'b101011100011111101001010;
rgb[15992] = 24'b101111110101000001011011;
rgb[15993] = 24'b110010000110100101110010;
rgb[15994] = 24'b110100011000001010001001;
rgb[15995] = 24'b110110101001101110100001;
rgb[15996] = 24'b111000111011010010111000;
rgb[15997] = 24'b111011001100110111010000;
rgb[15998] = 24'b111101011110011011100111;
rgb[15999] = 24'b111111111111111111111111;
rgb[16000] = 24'b000000000000000000000000;
rgb[16001] = 24'b000110100000011100001001;
rgb[16002] = 24'b001101000000111100010011;
rgb[16003] = 24'b010011100001011100011100;
rgb[16004] = 24'b011010000001111100100110;
rgb[16005] = 24'b100000100010011100110000;
rgb[16006] = 24'b100111000010111100111001;
rgb[16007] = 24'b101101100011011101000011;
rgb[16008] = 24'b110001110100100001010100;
rgb[16009] = 24'b110011110110001001101100;
rgb[16010] = 24'b110101110111110010000101;
rgb[16011] = 24'b110111111001011010011101;
rgb[16012] = 24'b111001111011000010110101;
rgb[16013] = 24'b111011111100101011001110;
rgb[16014] = 24'b111101111110010011100110;
rgb[16015] = 24'b111111101111111111111111;
rgb[16016] = 24'b000000000000000000000000;
rgb[16017] = 24'b000110110000011000001000;
rgb[16018] = 24'b001101100000110100010001;
rgb[16019] = 24'b010100010001010000011010;
rgb[16020] = 24'b011011000001101100100010;
rgb[16021] = 24'b100010000010000100101011;
rgb[16022] = 24'b101000110010100000110100;
rgb[16023] = 24'b101111100010111100111101;
rgb[16024] = 24'b110011110100000001001110;
rgb[16025] = 24'b110101100101101101100111;
rgb[16026] = 24'b110111010111011010000000;
rgb[16027] = 24'b111000111001001010011001;
rgb[16028] = 24'b111010101010110110110011;
rgb[16029] = 24'b111100011100100011001100;
rgb[16030] = 24'b111110001110001111100101;
rgb[16031] = 24'b111111111111111111111111;
rgb[16032] = 24'b000000000000000000000000;
rgb[16033] = 24'b000111000000010100000111;
rgb[16034] = 24'b001110000000101100001111;
rgb[16035] = 24'b010101010001000100010111;
rgb[16036] = 24'b011100010001011000011111;
rgb[16037] = 24'b100011010001110000100111;
rgb[16038] = 24'b101010100010001000101110;
rgb[16039] = 24'b110001100010011100110110;
rgb[16040] = 24'b110101110011100001000111;
rgb[16041] = 24'b110111010101010001100001;
rgb[16042] = 24'b111000100111000101111100;
rgb[16043] = 24'b111010001000110110010110;
rgb[16044] = 24'b111011101010101010110000;
rgb[16045] = 24'b111100111100011011001010;
rgb[16046] = 24'b111110011110001011100100;
rgb[16047] = 24'b111111101111111111111111;
rgb[16048] = 24'b000000000000000000000000;
rgb[16049] = 24'b000111010000010000000110;
rgb[16050] = 24'b001110100000100100001101;
rgb[16051] = 24'b010110000000110100010100;
rgb[16052] = 24'b011101010001001000011011;
rgb[16053] = 24'b100100110001011000100010;
rgb[16054] = 24'b101100000001101100101001;
rgb[16055] = 24'b110011100001111100110000;
rgb[16056] = 24'b110111110011000001000001;
rgb[16057] = 24'b111000110100111001011100;
rgb[16058] = 24'b111010000110101101110111;
rgb[16059] = 24'b111011001000100110010010;
rgb[16060] = 24'b111100011010011010101101;
rgb[16061] = 24'b111101011100010011001000;
rgb[16062] = 24'b111110101110000111100011;
rgb[16063] = 24'b111111111111111111111111;
rgb[16064] = 24'b000000000000000000000000;
rgb[16065] = 24'b000111100000001100000101;
rgb[16066] = 24'b001111010000011000001011;
rgb[16067] = 24'b010110110000101000010001;
rgb[16068] = 24'b011110100000110100010111;
rgb[16069] = 24'b100110010001000000011101;
rgb[16070] = 24'b101101110001010000100011;
rgb[16071] = 24'b110101100001011100101001;
rgb[16072] = 24'b111001110010100000111010;
rgb[16073] = 24'b111010100100011101010110;
rgb[16074] = 24'b111011100110010101110010;
rgb[16075] = 24'b111100011000010010001110;
rgb[16076] = 24'b111101001010001110101010;
rgb[16077] = 24'b111110001100000111000110;
rgb[16078] = 24'b111110111110000011100010;
rgb[16079] = 24'b111111111111111111111111;
rgb[16080] = 24'b000000000000000000000000;
rgb[16081] = 24'b000111110000001000000101;
rgb[16082] = 24'b001111110000010000001010;
rgb[16083] = 24'b010111110000011000001111;
rgb[16084] = 24'b011111100000100100010100;
rgb[16085] = 24'b100111100000101100011001;
rgb[16086] = 24'b101111100000110100011110;
rgb[16087] = 24'b110111100000111100100011;
rgb[16088] = 24'b111011110010000000110100;
rgb[16089] = 24'b111100010100000001010001;
rgb[16090] = 24'b111100110110000001101110;
rgb[16091] = 24'b111101011000000010001011;
rgb[16092] = 24'b111110001001111110101000;
rgb[16093] = 24'b111110101011111111000101;
rgb[16094] = 24'b111111001101111111100010;
rgb[16095] = 24'b111111111111111111111111;
rgb[16096] = 24'b000000000000000000000000;
rgb[16097] = 24'b001000000000000100000100;
rgb[16098] = 24'b010000010000001000001000;
rgb[16099] = 24'b011000100000001100001100;
rgb[16100] = 24'b100000110000010000010000;
rgb[16101] = 24'b101001000000010100010100;
rgb[16102] = 24'b110001010000011000011000;
rgb[16103] = 24'b111001100000011100011101;
rgb[16104] = 24'b111101110001100000101110;
rgb[16105] = 24'b111110000011100101001011;
rgb[16106] = 24'b111110010101101001101001;
rgb[16107] = 24'b111110100111101110000111;
rgb[16108] = 24'b111110111001110010100101;
rgb[16109] = 24'b111111001011110111000011;
rgb[16110] = 24'b111111011101111011100001;
rgb[16111] = 24'b111111111111111111111111;
rgb[16112] = 24'b000000000000000000000000;
rgb[16113] = 24'b001000100000000000000011;
rgb[16114] = 24'b010001000000000000000110;
rgb[16115] = 24'b011001100000000000001001;
rgb[16116] = 24'b100010000000000000001100;
rgb[16117] = 24'b101010100000000000010000;
rgb[16118] = 24'b110011000000000000010011;
rgb[16119] = 24'b111011100000000000010110;
rgb[16120] = 24'b111111100001000100100111;
rgb[16121] = 24'b111111110011001001000110;
rgb[16122] = 24'b111111100101010101100101;
rgb[16123] = 24'b111111110111011010000011;
rgb[16124] = 24'b111111111001100110100010;
rgb[16125] = 24'b111111111011101111000001;
rgb[16126] = 24'b111111111101110111100000;
rgb[16127] = 24'b111111111111111111111111;
rgb[16128] = 24'b000000000000000000000000;
rgb[16129] = 24'b000100010001000100010001;
rgb[16130] = 24'b001000100010001000100010;
rgb[16131] = 24'b001100110011001100110011;
rgb[16132] = 24'b010001000100010001000100;
rgb[16133] = 24'b010101010101010101010101;
rgb[16134] = 24'b011001100110011001100110;
rgb[16135] = 24'b011101110111011101110111;
rgb[16136] = 24'b100010001000100010001000;
rgb[16137] = 24'b100110011001100110011001;
rgb[16138] = 24'b101010101010101010101010;
rgb[16139] = 24'b101110111011101110111011;
rgb[16140] = 24'b110011001100110011001100;
rgb[16141] = 24'b110111011101110111011101;
rgb[16142] = 24'b111011101110111011101110;
rgb[16143] = 24'b111111111111111111111111;
rgb[16144] = 24'b000000000000000000000000;
rgb[16145] = 24'b000100100000111100001111;
rgb[16146] = 24'b001001000001111100011111;
rgb[16147] = 24'b001101100010111100101111;
rgb[16148] = 24'b010010000011111100111111;
rgb[16149] = 24'b010110100100111101001111;
rgb[16150] = 24'b011011000101111101011111;
rgb[16151] = 24'b011111100110111101101111;
rgb[16152] = 24'b100011111000000010000000;
rgb[16153] = 24'b100111111001001010010010;
rgb[16154] = 24'b101011111010010010100100;
rgb[16155] = 24'b101111111011011010110110;
rgb[16156] = 24'b110011111100100011001000;
rgb[16157] = 24'b110111111101101011011010;
rgb[16158] = 24'b111011111110110011101100;
rgb[16159] = 24'b111111111111111111111111;
rgb[16160] = 24'b000000000000000000000000;
rgb[16161] = 24'b000100110000111000001110;
rgb[16162] = 24'b001001100001110100011101;
rgb[16163] = 24'b001110010010110000101100;
rgb[16164] = 24'b010011010011101000111010;
rgb[16165] = 24'b011000000100100101001001;
rgb[16166] = 24'b011100110101100001011000;
rgb[16167] = 24'b100001100110011101100111;
rgb[16168] = 24'b100101110111100001111000;
rgb[16169] = 24'b101001101000101110001011;
rgb[16170] = 24'b101101011001111010011110;
rgb[16171] = 24'b110001001011000110110001;
rgb[16172] = 24'b110100101100010111000101;
rgb[16173] = 24'b111000011101100011011000;
rgb[16174] = 24'b111100001110101111101011;
rgb[16175] = 24'b111111111111111111111111;
rgb[16176] = 24'b000000000000000000000000;
rgb[16177] = 24'b000101000000110100001101;
rgb[16178] = 24'b001010000001101100011011;
rgb[16179] = 24'b001111010010100000101000;
rgb[16180] = 24'b010100010011011000110110;
rgb[16181] = 24'b011001010100010001000100;
rgb[16182] = 24'b011110100101000101010001;
rgb[16183] = 24'b100011100101111101011111;
rgb[16184] = 24'b100111110111000001110000;
rgb[16185] = 24'b101011011000010010000100;
rgb[16186] = 24'b101110111001100010011000;
rgb[16187] = 24'b110010001010110110101101;
rgb[16188] = 24'b110101101100000111000001;
rgb[16189] = 24'b111000111101011011010110;
rgb[16190] = 24'b111100011110101011101010;
rgb[16191] = 24'b111111111111111111111111;
rgb[16192] = 24'b000000000000000000000000;
rgb[16193] = 24'b000101010000110000001100;
rgb[16194] = 24'b001010110001100000011000;
rgb[16195] = 24'b010000000010010100100101;
rgb[16196] = 24'b010101100011000100110001;
rgb[16197] = 24'b011010110011111000111110;
rgb[16198] = 24'b100000010100101001001010;
rgb[16199] = 24'b100101100101011101010111;
rgb[16200] = 24'b101001110110100001101000;
rgb[16201] = 24'b101101000111110101111101;
rgb[16202] = 24'b110000001001001110010011;
rgb[16203] = 24'b110011011010100010101000;
rgb[16204] = 24'b110110011011111010111110;
rgb[16205] = 24'b111001101101001111010011;
rgb[16206] = 24'b111100101110100111101001;
rgb[16207] = 24'b111111111111111111111111;
rgb[16208] = 24'b000000000000000000000000;
rgb[16209] = 24'b000101100000101100001011;
rgb[16210] = 24'b001011010001011000010110;
rgb[16211] = 24'b010001000010001000100010;
rgb[16212] = 24'b010110100010110100101101;
rgb[16213] = 24'b011100010011100000111000;
rgb[16214] = 24'b100010000100010001000100;
rgb[16215] = 24'b100111100100111101001111;
rgb[16216] = 24'b101011110110000001100000;
rgb[16217] = 24'b101110110111011001110110;
rgb[16218] = 24'b110001101000110110001101;
rgb[16219] = 24'b110100011010010010100100;
rgb[16220] = 24'b110111011011101110111011;
rgb[16221] = 24'b111010001101000111010001;
rgb[16222] = 24'b111100111110100011101000;
rgb[16223] = 24'b111111111111111111111111;
rgb[16224] = 24'b000000000000000000000000;
rgb[16225] = 24'b000101110000101000001010;
rgb[16226] = 24'b001011110001010000010100;
rgb[16227] = 24'b010001110001111000011110;
rgb[16228] = 24'b010111110010100000101000;
rgb[16229] = 24'b011101100011001100110011;
rgb[16230] = 24'b100011100011110100111101;
rgb[16231] = 24'b101001100100011101000111;
rgb[16232] = 24'b101101110101100001011000;
rgb[16233] = 24'b110000010111000001110000;
rgb[16234] = 24'b110011001000011110000111;
rgb[16235] = 24'b110101101001111110011111;
rgb[16236] = 24'b111000001011011110110111;
rgb[16237] = 24'b111010101100111111001111;
rgb[16238] = 24'b111101001110011111100111;
rgb[16239] = 24'b111111101111111111111111;
rgb[16240] = 24'b000000000000000000000000;
rgb[16241] = 24'b000110000000100100001001;
rgb[16242] = 24'b001100010001001000010010;
rgb[16243] = 24'b010010100001101100011011;
rgb[16244] = 24'b011000110010010000100100;
rgb[16245] = 24'b011111000010110100101101;
rgb[16246] = 24'b100101010011011000110110;
rgb[16247] = 24'b101011100011111100111111;
rgb[16248] = 24'b101111110101000001010000;
rgb[16249] = 24'b110010000110100101101001;
rgb[16250] = 24'b110100011000001010000010;
rgb[16251] = 24'b110110101001101110011011;
rgb[16252] = 24'b111000111011010010110100;
rgb[16253] = 24'b111011001100110111001101;
rgb[16254] = 24'b111101011110011011100110;
rgb[16255] = 24'b111111111111111111111111;
rgb[16256] = 24'b000000000000000000000000;
rgb[16257] = 24'b000110100000011100000111;
rgb[16258] = 24'b001101000000111100001111;
rgb[16259] = 24'b010011100001011100010111;
rgb[16260] = 24'b011010000001111100011111;
rgb[16261] = 24'b100000100010011100100111;
rgb[16262] = 24'b100111000010111100101111;
rgb[16263] = 24'b101101100011011100110111;
rgb[16264] = 24'b110001110100100001001000;
rgb[16265] = 24'b110011110110001001100010;
rgb[16266] = 24'b110101110111110001111100;
rgb[16267] = 24'b110111111001011010010110;
rgb[16268] = 24'b111001111011000010110000;
rgb[16269] = 24'b111011111100101011001010;
rgb[16270] = 24'b111101111110010011100100;
rgb[16271] = 24'b111111101111111111111111;
rgb[16272] = 24'b000000000000000000000000;
rgb[16273] = 24'b000110110000011000000110;
rgb[16274] = 24'b001101100000110100001101;
rgb[16275] = 24'b010100010001010000010100;
rgb[16276] = 24'b011011000001101100011011;
rgb[16277] = 24'b100010000010000100100001;
rgb[16278] = 24'b101000110010100000101000;
rgb[16279] = 24'b101111100010111100101111;
rgb[16280] = 24'b110011110100000001000000;
rgb[16281] = 24'b110101100101101101011011;
rgb[16282] = 24'b110111010111011001110110;
rgb[16283] = 24'b111000111001001010010010;
rgb[16284] = 24'b111010101010110110101101;
rgb[16285] = 24'b111100011100100011001000;
rgb[16286] = 24'b111110001110001111100011;
rgb[16287] = 24'b111111111111111111111111;
rgb[16288] = 24'b000000000000000000000000;
rgb[16289] = 24'b000111000000010100000101;
rgb[16290] = 24'b001110000000101100001011;
rgb[16291] = 24'b010101010001000100010001;
rgb[16292] = 24'b011100010001011000010110;
rgb[16293] = 24'b100011010001110000011100;
rgb[16294] = 24'b101010100010001000100010;
rgb[16295] = 24'b110001100010011100100111;
rgb[16296] = 24'b110101110011100000111000;
rgb[16297] = 24'b110111010101010001010100;
rgb[16298] = 24'b111000100111000101110001;
rgb[16299] = 24'b111010001000110110001101;
rgb[16300] = 24'b111011101010101010101010;
rgb[16301] = 24'b111100111100011011000110;
rgb[16302] = 24'b111110011110001011100010;
rgb[16303] = 24'b111111101111111111111111;
rgb[16304] = 24'b000000000000000000000000;
rgb[16305] = 24'b000111010000010000000100;
rgb[16306] = 24'b001110100000100100001001;
rgb[16307] = 24'b010110000000110100001101;
rgb[16308] = 24'b011101010001001000010010;
rgb[16309] = 24'b100100110001011000010110;
rgb[16310] = 24'b101100000001101100011011;
rgb[16311] = 24'b110011100001111100011111;
rgb[16312] = 24'b110111110011000000110000;
rgb[16313] = 24'b111000110100111001001110;
rgb[16314] = 24'b111010000110101101101011;
rgb[16315] = 24'b111011001000100110001001;
rgb[16316] = 24'b111100011010011010100110;
rgb[16317] = 24'b111101011100010011000100;
rgb[16318] = 24'b111110101110000111100001;
rgb[16319] = 24'b111111111111111111111111;
rgb[16320] = 24'b000000000000000000000000;
rgb[16321] = 24'b000111100000001100000011;
rgb[16322] = 24'b001111010000011000000110;
rgb[16323] = 24'b010110110000101000001010;
rgb[16324] = 24'b011110100000110100001101;
rgb[16325] = 24'b100110010001000000010000;
rgb[16326] = 24'b101101110001010000010100;
rgb[16327] = 24'b110101100001011100010111;
rgb[16328] = 24'b111001110010100000101000;
rgb[16329] = 24'b111010100100011101000111;
rgb[16330] = 24'b111011100110010101100101;
rgb[16331] = 24'b111100011000010010000100;
rgb[16332] = 24'b111101001010001110100011;
rgb[16333] = 24'b111110001100000111000001;
rgb[16334] = 24'b111110111110000011100000;
rgb[16335] = 24'b111111111111111111111111;
rgb[16336] = 24'b000000000000000000000000;
rgb[16337] = 24'b000111110000001000000010;
rgb[16338] = 24'b001111110000010000000100;
rgb[16339] = 24'b010111110000011000000110;
rgb[16340] = 24'b011111100000100100001001;
rgb[16341] = 24'b100111100000101100001011;
rgb[16342] = 24'b101111100000110100001101;
rgb[16343] = 24'b110111100000111100001111;
rgb[16344] = 24'b111011110010000000100000;
rgb[16345] = 24'b111100010100000001000000;
rgb[16346] = 24'b111100110110000001100000;
rgb[16347] = 24'b111101011000000010000000;
rgb[16348] = 24'b111110001001111110011111;
rgb[16349] = 24'b111110101011111110111111;
rgb[16350] = 24'b111111001101111111011111;
rgb[16351] = 24'b111111111111111111111111;
rgb[16352] = 24'b000000000000000000000000;
rgb[16353] = 24'b001000000000000100000001;
rgb[16354] = 24'b010000010000001000000010;
rgb[16355] = 24'b011000100000001100000011;
rgb[16356] = 24'b100000110000010000000100;
rgb[16357] = 24'b101001000000010100000101;
rgb[16358] = 24'b110001010000011000000110;
rgb[16359] = 24'b111001100000011100000111;
rgb[16360] = 24'b111101110001100000011000;
rgb[16361] = 24'b111110000011100100111001;
rgb[16362] = 24'b111110010101101001011010;
rgb[16363] = 24'b111110100111101101111011;
rgb[16364] = 24'b111110111001110010011100;
rgb[16365] = 24'b111111001011110110111101;
rgb[16366] = 24'b111111011101111011011110;
rgb[16367] = 24'b111111111111111111111111;
rgb[16368] = 24'b000000000000000000000000;
rgb[16369] = 24'b001000100000000000000000;
rgb[16370] = 24'b010001000000000000000000;
rgb[16371] = 24'b011001100000000000000000;
rgb[16372] = 24'b100010000000000000000000;
rgb[16373] = 24'b101010100000000000000000;
rgb[16374] = 24'b110011000000000000000000;
rgb[16375] = 24'b111011100000000000000000;
rgb[16376] = 24'b111111100001000100010001;
rgb[16377] = 24'b111111110011001000110010;
rgb[16378] = 24'b111111100101010101010101;
rgb[16379] = 24'b111111110111011001110110;
rgb[16380] = 24'b111111111001100110011001;
rgb[16381] = 24'b111111111011101110111011;
rgb[16382] = 24'b111111111101110111011101;
rgb[16383] = 24'b111111111111111111111111;

    end

endmodule