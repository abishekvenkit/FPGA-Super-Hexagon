module audio_output(input  logic Clk,
                    input  logic Reset_h,
                    input  logic data_over,
                    input  logic audio_operation,
                    output logic [15:0] LDATA,
                    output logic [15:0] RDATA);

    reg [255:0] music [0:8355];
    logic [17:0] sample_num;
    logic [255:0] data_row;
    logic [15:0] curr_sample;

    // assign LDATA = curr_sample;
    // assign RDATA = curr_sample;

    always_ff @ (negedge data_over) begin
        if(Reset_h) begin
            sample_num <= 18'd0;
            // data_row <= 256'd0;
        end
        else begin
            // data_row <= music[sample_num[17:4]];
            if(audio_operation) sample_num <= sample_num + 18'd1;
            if(sample_num > 18'd133679) sample_num <= 0;
        end
    end

    assign LDATA = (sample_num[5])? 16'sd32000 : -16'sd32000;
    assign RDATA = (sample_num[5])? 16'sd32000 : -16'sd32000;

    // always_comb begin
    //     case(sample_num[3:0])
    //         4'd0 : curr_sample =  data_row[255:240];
    //         4'd1 : curr_sample =  data_row[239:224];
    //         4'd2 : curr_sample =  data_row[223:208];
    //         4'd3 : curr_sample =  data_row[207:192];
    //         4'd4 : curr_sample =  data_row[191:176];
    //         4'd5 : curr_sample =  data_row[175:160];
    //         4'd6 : curr_sample =  data_row[159:144];
    //         4'd7 : curr_sample =  data_row[143:128];
    //         4'd8 : curr_sample =  data_row[127:112];
    //         4'd9 : curr_sample =  data_row[111:96];
    //         4'd10 : curr_sample = data_row[95:80];
    //         4'd11 : curr_sample = data_row[79:64];
    //         4'd12 : curr_sample = data_row[63:48];
    //         4'd13 : curr_sample = data_row[47:32];
    //         4'd14 : curr_sample = data_row[31:16];
    //         4'd15 : curr_sample = data_row[15:0];
    //         default : curr_sample =  data_row[255:240];
    //     endcase
    // end

//     initial begin
// music[0] = 256'hc2070e07f703f4ff36ff1f00b400c100d3004700d4fd21fcaafb73fb27fbe7f9;
// music[1] = 256'h00fa4ef79ff41900670ce00a9c09220a7207b6067805e503c7034d025801a800;
// music[2] = 256'h83ffe1fee0fdbefd50fde5fb6afb6cfa82f901f98af764f643f582f430f4f4f2;
// music[3] = 256'h3ef2b4f11ef10ef1e2ef16eff9ee3ceecdedc3ec01ec00ec20ebcbea54ea7fe9;
// music[4] = 256'h49e99be8d2e8f9e7e8e6f7e86ae2bed33bcff1d09ecf3acfaece07ceb9ce6bce;
// music[5] = 256'ha9cedece02cefbcd4ecdf3ccf6cde7cdfbcd7ece31ce00ce78cd4ecdfecddacd;
// music[6] = 256'hb6cd2ace65ce9aced0cedacef5cec1cf50d0d8cf5ad01ad1dad07dd153d287d2;
// music[7] = 256'hfed23cd37ed3dfd30ed454d473d4ced47ed5d4d565d676d8e1daf2da88da68db;
// music[8] = 256'h37db36db4bdc9bdc7bddb7dfebe142e20de237e3fbe232e364e410e36de3dbe3;
// music[9] = 256'h84e3bee5e0e236e753fd2309c5051906b8063c064d070008120ac10a4d0a040b;
// music[10] = 256'hbf0ad80a1f0bb20aa40acb0bbf0fe7118a109910a010761075117911cf116f12;
// music[11] = 256'h8f12f3129012b41276132d13241369139d134d1405156a1597151d16a116af16;
// music[12] = 256'hcb16e11603171f17f816191779173a17db15a5153617b11763184919b4179516;
// music[13] = 256'he516c8160a17a2175a180618a5155f147a15ec14f2114611a711cb109f11ce10;
// music[14] = 256'h9a124b1e0126fe2425251425922447247a23f223b923a4244c24522372272e1e;
// music[15] = 256'h7908530349065e04ae05410692055b06860574059d054605ba0589059f05a805;
// music[16] = 256'had053b06de05e005010686062108020888073207220668061706b40527066005;
// music[17] = 256'hf5055006530694072a003af45cf2b4f3e8f1aff148f180f018f1c0f016f052f0;
// music[18] = 256'h1bf047efe1ee00eff4ee52efe8efecef7af178f3ebf23bf2d7f18cf085f0fbf0;
// music[19] = 256'hb1f08cf027f03af076f017f07bf0a1f01af043f035f0f4effdefe8efe3efabef;
// music[20] = 256'haaeffaef26f0a0f0b9f034f010f0f3eff8efa4f00ef1f0f0ebf0e0f0def071f1;
// music[21] = 256'h06f215f2fdf113f27ff2a9f2a7f204f3d4f2eef2cef313f474f4cdf4f1f470f5;
// music[22] = 256'h1bf572f57df6fdf596f569f5e8f5e2f750f822f8adf89ff8cff866f814f88ef8;
// music[23] = 256'h3af7c6f5caf531f716fae9fa9afb70fe9dfee0fd40fec2fd94fe76ff3dff89ff;
// music[24] = 256'h08ffcafe20ff37ff9eff04fe48fc50fd27fe43fe08fe5dfdebfd85fea7fe2aff;
// music[25] = 256'h82ff90004401c800350051fefefd3e00a7ffc5fd36fd33fd77fe8cfe8cfdfffd;
// music[26] = 256'ha6fe0affd8feb5fe55ffeeff54001cfe86fbfdfb64fb7dfa69fa48f946fadefa;
// music[27] = 256'hb6f9d3fa4dfb7dfbf4fb93faa4fac1fa00fbb9fca2fcfbfda8fe2bfd51fcfef7;
// music[28] = 256'hf5fed0148d1d221a25194119dc1b2f1a1a14f1155f1cbf1f011e2b19e7163c14;
// music[29] = 256'hda0ff30c2d0a3f0c7f1329152d0e95026dfb98ff7f055f01ddf436f03800fe14;
// music[30] = 256'hc41b261aa11a7a21d326e11b000d4c10a818d412d600b8e988e278f88211801c;
// music[31] = 256'h34200a1c9d17ff16630cc9fdc9f98bfb02fc3dfbadff7e0a0511670d7407f70d;
// music[32] = 256'h6a1bc61b2311a1061107a916e2207118990482f196ee0cff231c273b0149013f;
// music[33] = 256'hec28fb168e159024bb3a37471b39d51d2e0f8e0dcf12051ba920fa26892c272e;
// music[34] = 256'he5320e37c62e46233924062cc32e4d28891edc2192349740393744279e1e3a1b;
// music[35] = 256'h701ede21f71f69219c25a42ad12f692b7c1cf810cf109813d5178b25ff379346;
// music[36] = 256'h5d4e834cce41d73c6948585a4b667363ca50373ab628541e3614f10245ebeed3;
// music[37] = 256'h31cd4fd255ccb8ca63deb6eea1f0ede656d189c42ac537c8f4cea0d365d82ce0;
// music[38] = 256'ha1e623ef7cf86102600cbc171f1bee092e04f2121e1d5b28073147360f3fa53f;
// music[39] = 256'h043af22b3b1df21efc1c8c11270b79056e027b031904970411ffeef744fbeb03;
// music[40] = 256'h8507fa0075f992fe5507970f181c1c21dc1af40bb5fc9e079122ac295d28812b;
// music[41] = 256'hc2216b171a26c148d466316e806467534846234604416833cf27a518fa0e3917;
// music[42] = 256'hf233f15af66d8769896607709e778d6fd6660d691b73cf7bae770375ac79757a;
// music[43] = 256'h9e7c7a7d7d7cf27dc579b172666fbe72277aa57885719670346da75b6b4c2a52;
// music[44] = 256'hff57634d6a41403b3f4656617e6bc768d96c346cef657b5b69510c5439598857;
// music[45] = 256'h185256501553234f1049ec484650b559f05572477338672e59289d1ef812ea06;
// music[46] = 256'h1804dc07effbc6f161fa58042306d5faa1efbbfb4e12a31c6519390e8e00f9f7;
// music[47] = 256'h56fcd00a74104205a7f9b8fa2dff32f796e8a4e532ed34f03fe983dec2d6f3d6;
// music[48] = 256'h0bdfa3eaf4f333f7b1f870f3c7e530de76d9c7da02e6a2e3c7d75fd6f8d355ca;
// music[49] = 256'h71d0aff0061094171d0dc408920fe50930feb5fca5fc48ffa70d31283d398531;
// music[50] = 256'hf32365178c0be70af516d82b323c2e401743394ae74d3b425b2a781f8827b42f;
// music[51] = 256'h9337483e77392c3101216c07e7022c1a57385a47fc39bb2552253132cb3a5634;
// music[52] = 256'h2f1f69106d177c25732a0824ba170313211f8f300234542e442b0a2dcb340535;
// music[53] = 256'h453187399f3e053c733c7c3a5936a1351933f02c562868230e1d3313e007cc08;
// music[54] = 256'h1a0c0608b7069609160e4a0af4002efc0ef6b8fa1309700b3705a8014202d003;
// music[55] = 256'h130341fecbfcdc03370fab23da2be21ceb17e71f5027b6261f1c0213d80af20d;
// music[56] = 256'h3c1335042100ac10611b4b18dcf84ccb2bc159dbcbebc9e0a0db2ef279071908;
// music[57] = 256'h670479068f08f3050e05900395ff62042e0362f3d4e6bbe130e58ce56ad4b2c2;
// music[58] = 256'haec7d9d992dc64d706d984db89e28ae305dc50d87ed293c910bfdebe2ecb48c4;
// music[59] = 256'h88aecca245a1f0a7e9b168bea7c373bcdac435d69cd4a2cbc6c754ca02ca53c3;
// music[60] = 256'hbcc59cc8a3c8e6cc79cc58cb8cc297b039ad3ab4bdb526b4cebfadd336d4a1cf;
// music[61] = 256'hc6d5abd486cee9cc96ccc5cc98d588e2fad508b75cacf4b70bcd61dbafd25ebf;
// music[62] = 256'hb0b5d8c133d68ddc25de4bdc09d7bdd582d005d089d67cd986d8cdd22ad569d7;
// music[63] = 256'h09c80fbc29c235d360dbd8cc28b64bab45bcf7d9e0e303deeacf6fbe18bc47cb;
// music[64] = 256'h82de56dbc2c212b76fb325b313bf7fc664c8f1c294baa8b961b864cc9ce6a7e6;
// music[65] = 256'h04ec81f9ff004c08810d5e127d12eb14d30f4af7d2ea01ed7aeed6efcaec61ec;
// music[66] = 256'hc1edccee2cf1e0effaf9ac0f23184d17681ab21ef516a1fd14f1be01b714a31d;
// music[67] = 256'h4322f8235420651c5e1d6f199c0ae9f5b5f55e108b1d591cd01adf177f1a9b14;
// music[68] = 256'hcb09cafd02df7ec8f7dc5d09df1b1410bb04c9fc25f986fe0606cefa51d7d1c5;
// music[69] = 256'h68da3afb570757f273d9e9d534df24e100e03aef9bff4dffe0fc8f071e107cfe;
// music[70] = 256'h8de52fdf92e0d3e0c1ec36073a17dc0c55ffaa030d0956fffef21eef04ee6beb;
// music[71] = 256'h7cf5250b1912630a3407b20a350511f5eef108f92cfadbf741f702f740eff3f2;
// music[72] = 256'h6c0edb1c460c9af291f00d0ba5204e1d52047aec6eefaf09b9227020670a6afb;
// music[73] = 256'hf4fa6908f2148a0ecef9d5e9bdee6803fe102d0906f7ccee1cf9780d13141107;
// music[74] = 256'hd1f2a7e5efee4c00520514033102f50238f475db03d200cfb9cf21d80bdaedd7;
// music[75] = 256'h66d5b6d0b3cecdcb6cc6c2c525cb7ecc34c740c2f6be91c079c4edc3b5c057bc;
// music[76] = 256'h75bc51bf27be08beb0bf07c2edc18fbf37c294c135c5d2d7d0de2cdb35e9adff;
// music[77] = 256'h7e05baf66be19bd901ec7604d708d8067d087c07cf07c1071007140378fb2dfc;
// music[78] = 256'he2fef7fd09ff7bfe65fcf4f76af4c1f745fa04fa8afabaf991f710f53af285ed;
// music[79] = 256'h3ae912e81ee84bea58ebf8eb20f0a4e2eac0cbab1da680a571acb0b219b28cb3;
// music[80] = 256'ha4c6b0dc1bdd6ddae9db41d637d009cf5cd849e448e638e418e1b6db8dd40fd3;
// music[81] = 256'h62d671d7d8dd33e603e8ffe3eedf40e434e620e2c4e133e5d5e909eaf2e95feb;
// music[82] = 256'h27de22c616be22d143ecfbf992fb01fedafae9e27fc751c500dc00ef31efd0ef;
// music[83] = 256'h49f2e0efe7f135f302f2c0f4bbfa62fff4fb2df42eef67f1caf8e6fafbf622f5;
// music[84] = 256'he4f83efc99fd24ff7cfeb7fea4fd3800290be301b9e312d921e3c9e688e628f4;
// music[85] = 256'h530b3b12a7ff2eeb76e671ed79f3e0f31aff0f0c7d09e8097f0d1d0fd517ea1a;
// music[86] = 256'hd91688178f1ae21cb11ef51d521c851c2f1cb21ec22266209d2071272c2b2c28;
// music[87] = 256'hba26b62a3a21400ad6ff670a80200c2a541b540af906a1078e0227048416372a;
// music[88] = 256'h8d33a730d121fb1b6a30b6498c4d6f464f482c4a7344dd40be420c4ae94c2849;
// music[89] = 256'hb84a8b4d7654d25b1e5828554455ca59d05e575d3861445c814d5b4a30414630;
// music[90] = 256'h1b32493efd3c073ed44e695fab667a58ba437d3d9e363b34a12de41a4810320b;
// music[91] = 256'h0717282942269624a926a3232821561d1a1e1920df1fce20082174227a24ce26;
// music[92] = 256'h6828c62762295b2ba3222e0d9e01330f8a26f43336353a386539cf26da0ed108;
// music[93] = 256'hb00d140e6210002195315830412de234ce33bf22a514501a7d30c43cbf35a830;
// music[94] = 256'hf9347a376a322a2db22f93324d33ad35f3337c30ac2c6f29842ee726690c8701;
// music[95] = 256'hce09fd0f300f9a142924cc254e15fc01def9db09e01f3624001438fe54fa5906;
// music[96] = 256'h5416311aaa08e2f769f11df0e5ef3af39b07671749149012440ed308b30b840f;
// music[97] = 256'hcf10790c670adb0ce60b540e34046ae501d8a8e94b046e0f50fbc4dc28d3a4da;
// music[98] = 256'h76e5e2ea1ae482dd7fde2fddf4dac4dcf8df2bde60d726d57fd3f7d325e56bf4;
// music[99] = 256'h1af59df446e8dbe1bffb2c103714ff162c11cf0dc10c2c0c590ffe0b910a9efe;
// music[100] = 256'he7e5e1de58e14be6c8ecc4ec55eb04e2ade53dfd910593073008d5fef4fa2bfa;
// music[101] = 256'hdcfe1c0378ff9c01f8fe2bfd25f98adf37d42edb1adea3db7ecba5c4e2c6eec7;
// music[102] = 256'h6edc3fead7e850ecd8eacee7cbe64fe953e783d045c47cd38ce4d2ef15f524f6;
// music[103] = 256'h6cf329e6c9d5d0d238e518f8f2f8e7f8b7fc5cfccdfbbcfd4d0228032004a604;
// music[104] = 256'hb8f3abe1ffe9fe016f0f240bd807520f0e0e92f9cde981f2eb08021500114c12;
// music[105] = 256'hbd1a0c130ffd7bf1e4f5acf604f5c000f3169623af14d2fde9f674fbe9fdb6fc;
// music[106] = 256'h400f032544233d22fa23ff1e1f1b871e8721740e79f945f994fbfbfa72ff6e0f;
// music[107] = 256'hd120ab1e4e0d8b00f7fef6fe6cfcca035a187f26f21e5d07b8f7ae040f18761a;
// music[108] = 256'h480c6cf5f0ed43f3a0f333f1ebf20b05de138a075fef97e582f6bb0a810e5f0c;
// music[109] = 256'hcd0f1014a70361ecfaea9bf9a509d30a1ff889e68ee060db9dde3af3700a511f;
// music[110] = 256'h151ea003c4f3c4e928e184e603ecfdea9ce4f7e151e6f0e92ff70b0bfc0ff8fb;
// music[111] = 256'h08e006d99fdecddf13e37fe774e6bbe4b2eefdfe97fff8edf4da4dd6f8d895d7;
// music[112] = 256'h19d9e7d906da8de12bf2b90420f6dfd263c8aec8bec3cbbcb1c00fd747e3fbe2;
// music[113] = 256'h33e55ce6bfe2ebde93e191d878c515c175c2babf4ec0d0ce0fe32ee8b9e469e8;
// music[114] = 256'h3aeb09d8f2bbafb680c044c41dc73fd6fae21de1bfe0efe581e27bcce6bb9fc2;
// music[115] = 256'h15c88fc7e6ce4fdf7cea58df14c8cabb91cb89e73ef326ef52e9f9e6abd83ac5;
// music[116] = 256'h86c5d5d509eb57ef84de25cb17c3edd18de54be7ded743c703cb4edd1cefc0ee;
// music[117] = 256'h15d73dc268c583dbe0eb84e61dd08ec00ccbb5dee7ec85e86cd36bc9eacb9ecf;
// music[118] = 256'h82cec6cb97c7dbbb08c47ae482f87bec10d0e2c2f7be7aba55c2a1cecbd381cf;
// music[119] = 256'hdbc6b0c234c57ccac0ca48cc08d0f3cc10c9eec4ffc0dcc5eacd24d024cd89cb;
// music[120] = 256'hf2cd38cd49c898cae2d7a9de4adc5dea15051e12990f6709310628fa6ce7d6e3;
// music[121] = 256'hb8e55bdd4ad696e7cd07a710770b92096b0168fbf5fa01fdc900a503b107e708;
// music[122] = 256'hf906d202a2fb5ff6c0f638fce8fd11fbc4f9dbfa9cfd09019bff34ef32e4f9ec;
// music[123] = 256'h4ee6c3ccf4be7bc59fd681e3e4e1d8cfbac134c9a6d841de63d38bc523c5c3d5;
// music[124] = 256'habe6cae2d8df6fea71ec3de88ce30edc55da4cdf7be324e9e6eeaaec5de970e8;
// music[125] = 256'ha8e50fe476e4d6e747eb42ed2aeb2fe386e2d1e292d5b3caedcd44d3b6d36bd3;
// music[126] = 256'h5bd20bd29bd256d35ed5c8d592d849d862d50bd30cca7bd748f4b3f4c0ed6ff0;
// music[127] = 256'hcef238f426f357f399f5f5f51ef26ef152f8a1fcbbfb4df8e0f5d7ef4cee0ff7;
// music[128] = 256'hf3f9bafb83f32fd926cb71d7caf35aff50f85ff5cbf12ff45dfa07fd16fd7cf7;
// music[129] = 256'h51f560f297f6c2fde7f15ae05ed6e9e019f534fcc40014ff4ef9a2fa69000e06;
// music[130] = 256'hd7040b0026f902fb6d05070bf61695235022da1d9722c621ca0d5b02ed05d506;
// music[131] = 256'h9401f1069d1f642bb2296526f61def1f311d7117af1a15200428011c99069401;
// music[132] = 256'h60020a032c01130de71de41d611eda20ee211b27e02a3d27ce1de81ae6136306;
// music[133] = 256'he706bc092e0691094e0911f9daeaaef0f5046c12a70ad1f408e26be8f0fdec02;
// music[134] = 256'hdf03950c761221144312641056038dec63e72bf6e3089b0af9f7cae735e697f6;
// music[135] = 256'h610b9011c911f412c113a313fa0e910b680ab80758050b06fb11701748025eed;
// music[136] = 256'haae59be2efe8d5f03cf170e869e04ae54fedd1fe6f15a1124504bd04b10c0d05;
// music[137] = 256'h70ef94ea3def05f054f458f328f023ec74e7b2e8a3ed2a030d166012230fd40d;
// music[138] = 256'h910efc125c122b0c6d06fc1126185f0491f150f2e2072b15500d1f0a7c0e5c14;
// music[139] = 256'h72188817d903c7df05d600ed8308010eb1f629dc85d25fe20dfd370b500ecc0d;
// music[140] = 256'hd50ca307c3072705f8f109ed83ff5a17ec28d82c602f9b336234373327340d2a;
// music[141] = 256'hdc104609ef14bc1acc1587155a21202306257c30a838bf37c822b4131012db0e;
// music[142] = 256'h4815fe13180b8705cc024b053002e60ec822e91ed3190a14ad0050e80bd88dd8;
// music[143] = 256'hdfd903d019cb8ae040fc4f049104b402adfa9ce8b0dc36eb0dfc1002c6fc77e9;
// music[144] = 256'h16dd88e6b2027416e20df1fa2bf15dfd64112417dc17ae19e41819148b122819;
// music[145] = 256'ha911e9fb17f79905a915cd19e70afcf64ff46b07c8209f25970f55f931fa760e;
// music[146] = 256'h2c1fec1cf20f8a0859082a0354fdf2fe45018201a2ff6902eb06d102220036fd;
// music[147] = 256'haffae7fa69fa3e0ebb257623b41ba91cad20051328fa49f765fd5dfd41fbb1f4;
// music[148] = 256'h46f33af884fa9ff985f756f814fb4ff9dcf921ff52ff4701ff03220b1722882a;
// music[149] = 256'h841f1220df28f12d502b4627a9281f2b232cdd271c24f124051732fa40fa9c24;
// music[150] = 256'hd146d6480436481a760eda1c1f352243cd459946ef435a3ee1378b38693de33d;
// music[151] = 256'hbc3d3a36d830df36ee3d1945c63c0325cc167c1fc232e7331f2e2d330137a934;
// music[152] = 256'hfe301835333ab43b5636511c4205e801e800dd002e0374002bfc89fca0fd29fb;
// music[153] = 256'hcff95e0ba7234320451bcb2368278a2b1627cd1b6d133d12a21fab28932dfb24;
// music[154] = 256'h1704a1ee09f43e021fff2dfb810ead1641158f18581558122f11e2101f09cbf7;
// music[155] = 256'h42f454042216a31964158713421352147618f61a6b0d95f78cf2e7033318861f;
// music[156] = 256'hdc24c525091f4c198a122511301330194b1cf208bbf66efbfe0fdc243525e90d;
// music[157] = 256'h0ff4bff88611be1e0121dd23692a1f1e0705f4fe130315041dfe2d0229141618;
// music[158] = 256'h4515a819601b2e0d33f61bf01df462f5eef9800c711fa11d7e1cc4212f1ef417;
// music[159] = 256'h28157d15a10851f81afea50b8e0b7802d4026303bbfb65f928f9810764211d29;
// music[160] = 256'hda1c4e05bbfa930aa421652e4923740a01004d0dbc203b23491395fccef4b701;
// music[161] = 256'h940f9412ae0259eacae7adfe94121c11bf0920fd50e417d0c6c0cabf55d344df;
// music[162] = 256'h8de36be68de56be749e271db0dd16cbaa3b059b04aae91b3e6b4b2b2b2afd1a7;
// music[163] = 256'h14a513a695a9b4ae09ade4aa8bac56ad62ace7a95da53ba14ca37aa6aba4b3a1;
// music[164] = 256'hc2a411b7e7c897c5bfb608a7ada157a5c3a4abaf61c3dec722c328c320cc59cd;
// music[165] = 256'h45bafeabb1b02fbbfbc395cdd1d6a6d979d385c654c1b5cb0bd7e5d825d064c3;
// music[166] = 256'h67c092c9a5d356d592d36ad671d94cd401cd19c823bdb6b4bab58bb0d3a835b3;
// music[167] = 256'h31cec5dff3d61ec0d7b313bbcdcc46dc47d957c8dbbf1abedcb950b2e0bb60d9;
// music[168] = 256'h9ee2e6df29e44be00edbb9d620e1fdf99f024e049704a6033109c207c002eefc;
// music[169] = 256'h9dfba1088c0954f26cdac4d6b3e967030a0a53f8eae759dea2d8e5dd1de5a3ea;
// music[170] = 256'hd2e79de217e7c4e649eee903d30a48fc26e737e4efef02f7b1fb9df987f580f5;
// music[171] = 256'hf6f4b7f66ff537ef5eec20f20efbc8018105e6fd70fcd40153f21ae30be0dfdb;
// music[172] = 256'h26dcb9dfafe6d6e5aee309f7b80675096e0cad0b3c0b98073c0478fbd7e320db;
// music[173] = 256'h67e165e329e2cdde1ce101e19eeab6022a053c02b0042efccdf821fbd701d506;
// music[174] = 256'h97066f0adb098a0ba2036de46dd263dcabf2e7fd64fa7bfd17069a0162e70cd0;
// music[175] = 256'h63d749f42b0cbc0c3f06f102d6f507e2ccd81ae69ef9ac0029fd5cfc84019cf6;
// music[176] = 256'h22e42be171ef4f02670392018204f7031a06a701d7fbf4f9ee00c90a0af88ee0;
// music[177] = 256'h7ddb12df6de001db75f02e132a138cfd29ef60f058f15fee52f5ba08f7173b0a;
// music[178] = 256'h03f2dcebd8efbcefb9e86def1406b6118107d0f511edbfeaaee5e0e370f4f106;
// music[179] = 256'had08590ed71622185213b10d4a0abcee61d3e9dcb8efb7fb7ff29ed84cd17cda;
// music[180] = 256'ha0dfe9dac0dcb1ec37f7bbeee4dcffd610d9c0d598cfa7d2b6ebc302a3fc5ce7;
// music[181] = 256'hadd750d10dd0f2d211e17cfaf90436f43bdf7fd619e08eeffdf7dcfdb00075fb;
// music[182] = 256'h18e5d3cf86d206dbeddeabdcded408cddcce73e6e7f95df419e43dd771d633d5;
// music[183] = 256'h5fd3bcdf2ff3fbff41fb63eb32e3a8e104dc89d79adfa3f1950085fb0dee0eec;
// music[184] = 256'hbbe864e1d9dde4df64e3b0e280f07705de07eaf9c3e10fdc8ff3d60562067301;
// music[185] = 256'h2004d7049ef334e3acdf6be060e250e9bcfa160791fa5fe47ddaebde02f11605;
// music[186] = 256'hb411a823c02a221682035900720354ffcbf66305081d0826d527782803295618;
// music[187] = 256'h7dff17f8f7f6dff95e026208a006eafd4c0594181e1e5513bd026ffd0d094b17;
// music[188] = 256'hcf0b86ed0fe6e1eb1ae728dfabe2cefac10dbd0570f266e4ecde4fdef4e2b9f0;
// music[189] = 256'h6703cd0812f983e62be133f28909020b2ef97be39be0b4f0fefcfd066c0bce0e;
// music[190] = 256'h2a10bcf82ae564e6e4e481e6f2e870e9ceeb60e7a8e330df65e0b0f3c3ff92f9;
// music[191] = 256'h0eeaaedb4adac3d74ad500e70b00ef07a5f8d8dfb8d367d689d831dc53e687ee;
// music[192] = 256'h98f3a2f30cee19ea0deb6ced44efe0ff1a1997207a15ad033a02ed127615530d;
// music[193] = 256'h2e15e72425254a208320df196410f90ce60d4c057df415f6e908ef16ec0b11f6;
// music[194] = 256'h1bed5ee666e2a5e134f4da1b0e29e628892c762b1630a92f0e31c130382d8231;
// music[195] = 256'h5a25931acb1efc1e5d1fd51a9719001fb72b3045e34ee747d949aa524d50753b;
// music[196] = 256'h7d2de137d24b3756554fa735a31b4f1d922941292b2e313874342d2808209b23;
// music[197] = 256'h46381b47023e1235b4396141ef46ce494645ee31461e7e21d03796466942e23d;
// music[198] = 256'hfa44ae473b3614221521de2f1a435541f92ac2213028e32d692bf925af238021;
// music[199] = 256'h6128123a8c46da40ee30bc29b125301a38116813c5153715df224e342a36ed2f;
// music[200] = 256'hab2d322c7a166afa44f8e001f907860f831d442cd622380959008c036a0266fe;
// music[201] = 256'h7fffa2035200e903e6143c1a7215ce172c1d79151dff19f59dfc49ff30fb3c02;
// music[202] = 256'ha615db1c5e193e1bcc19f7094cf0ecf323186f2eb732ee2731168b1847271f33;
// music[203] = 256'hc22d6f1a9210b30ef90b84039305fb200a35b333aa30ff31f62bf716320a8013;
// music[204] = 256'ha1253334e12e521b2311a814bb1f8f1e2107b8f32cf3affd700b210caef95aea;
// music[205] = 256'h12eed0f6e3f8f2f6d5f1c5ef0eefe6ea9ceb02f0e8f3adf107efb4ff50127610;
// music[206] = 256'h03ff8aeb59eec7051f1ada181d03b4f517f4f0f2f7f78dfd57ff6aff5ffe74fd;
// music[207] = 256'hf8fd3f015502be002d01b603d605660678040401060bc01b9d1e4a1ea01cca17;
// music[208] = 256'h6a18b11c5c22f820191e741732fdfaed78f748ff40ffaffb90fb42fc36f9dffa;
// music[209] = 256'h7cfd37042d1115131912ad19881c251abd12f009310c3d13e518a7188413b711;
// music[210] = 256'h930dbe0fd215b50cd7f87eeb7500d1275e306e2ac530fe2fd424022512258013;
// music[211] = 256'h9affccf875064f172a190f1bb21de61c4a1bca1af116a402ddf32afe2011da1b;
// music[212] = 256'h2d1a9d188c17a0144814b00c87fb3ef072f385f25cec10eb2ede33d02dcff2cb;
// music[213] = 256'habbd8db2b0c15bd655d710d312d709d75cc30bb21ab3c0b4d2aee0afaec53cd5;
// music[214] = 256'h68d282d14ad470ceb1b8c8aa95aa82a5d4a85dbbf3d63de3dcda5ed7d9d55ed8;
// music[215] = 256'h86de13de0adc31d867d7e8cdddbbd5b764c344d349d421c61abb53c03ed460e0;
// music[216] = 256'hf5db6bc634b301ba79cfbde082dbf5c835bf58c04ccd50d725d429c5cdb79dc0;
// music[217] = 256'h15d48fdfedd873c071ad46bc1ee086ee5dedd8ecf4eb1dedece9fce986e0bbcc;
// music[218] = 256'ha3c6dac519d53ded4cf1c3ef82ec80e777eaf8f02df205ee7cea41e736e80bef;
// music[219] = 256'h34f617f9def368ef00ed99ea4ceebcf73cff6e0143fefbf018e801ee22f7ccff;
// music[220] = 256'h60f552e55fef0efd4701c404bb010df1addc93dc4cecbff79af6e6f146f40cf8;
// music[221] = 256'h8efe8a062a0a6c0945011afbabfb42fdd1fd10ff01040008c00878057ffe9cf8;
// music[222] = 256'h6af6d2fc2704e805a20877071f01defd0aff3f0324ffebeac4e366f7ee07300a;
// music[223] = 256'h95fb3ce439dfe8e319e49de750f76f075d0233f954f72af737fcc0fa8df94ffc;
// music[224] = 256'h46fa4bfbc1fa4cfb5dff04009502ab0149fea3f93ef1dbf1f0f75ef74bf321f4;
// music[225] = 256'haef5d1f431fcd1f7dbdfc4d53ed61bd4d0d325cf8ed33bea8002a815e31414fa;
// music[226] = 256'h75e4c0e639fcbc11a313ee0fd01027110f141112b8096b0aa816481f4a1d0216;
// music[227] = 256'hd60a08055d099e13371e6f1c0d15ec0973f561ed3df38ff718ef41d941d044da;
// music[228] = 256'h26e9c8f179f1ccf9f9fe10eb6fd230c9d1cb08ce13ce40d30dd4d1d474e61af7;
// music[229] = 256'h4ef723efc8e619ea0af3d9f36af1acf1f9f38af449f2e4ee83ee0ef178f202f9;
// music[230] = 256'ha2fd1dfc89f6eaec0cf2bff0d9d954d19bd651deb9e281e876fbbbfde1ed20e1;
// music[231] = 256'h45df39f4120579fe1df44bf306f9f8f1f0e108e27df3e9012b01d1fbc1fa76f9;
// music[232] = 256'hb9f767f664f448f81e02e104380000fb53f960f9f1f7e4f6d6f3f7f3d1edceda;
// music[233] = 256'h11e0befa5c0d9116df08eaee2ce8c7eeb8f1c4f041f421fa69fea009db16ee0d;
// music[234] = 256'h19f3afe5bceb57f6b8f7f6f661068911f20c7a0c6c0e3511b51063066201bcff;
// music[235] = 256'h86fb96fb08fc56fce9f97ef9e60189f9cede94d1acd410db95df47e444e443dc;
// music[236] = 256'h1de238f534fba6f549f6d4fbbcf2fede62d79ad858d852dbd3e95dfc4cfc9ee7;
// music[237] = 256'h0dd67cdc64f4e4048605e3007bfc87f679f5ebf7ebf590fab703aa052506f403;
// music[238] = 256'h42f952e419d403e24cfeb70bcd0dc6103112130454ea43dfb3ec5e008b040df6;
// music[239] = 256'he8e374e288f4c4044a05aff992ec4be81ae6b3e031e345e930e698e404f27a01;
// music[240] = 256'h85028f02f3119822a828ee286325d329e7320c24c1062cf91efb46ffd9022e13;
// music[241] = 256'hc02a472d97158efcc2fddf0b840abc017efcc0fff4087b0b370bb8040cf244e5;
// music[242] = 256'hc8ee0d0a7b1c6e170d0a4c03780286f82be687e514f658fd53ff630a2d11f110;
// music[243] = 256'h6e14a6145c08f7f2bce9fff79e0b6b139f0592ee73ed60fe52063405800d7819;
// music[244] = 256'h3b1a261b8e24992d8d314231232639136f1430206d17db0c6313fb2595378534;
// music[245] = 256'h8f20e60ef709220889fee7ff31147e24d323351d9816c60842faa6f66efa65f6;
// music[246] = 256'h21e930e7a2ea98eaaff99b10211c381664039ffd2e0c381d8f23a31f95216f24;
// music[247] = 256'hc724fb37db471d3b652ddd2a66272324d225ac27b624c82b9c475f5f6f5a6540;
// music[248] = 256'h0428ea2845421f54564c4334e925c435904f6358ac53654d5842452df31b2819;
// music[249] = 256'hc71f26247a215120351b2f1679244037c63856341f3b8a404f31b6188e0eb61c;
// music[250] = 256'h732da22f8934f93e133e482b4c16fb0d89077f076710e510600f340ff00c020d;
// music[251] = 256'h9a0a23078306ea118c29503263275217100f5d182526a22a2424f821cc29f723;
// music[252] = 256'h1d15980ee4133521e91f66126a0825048203e3fea203a0171226c622090ee4fa;
// music[253] = 256'h9efd1e147526cb2757262f28fc2ad329a425f723e41db41c701f6419a5177619;
// music[254] = 256'h32176f166817b517ec16781ff6309d350729621c0e180816ef11320ee40c900b;
// music[255] = 256'he10d131c6f3045361326a31a9c186107c6f4c2ed56ea6decb6f7e70f8c1d8612;
// music[256] = 256'hff0ae00a800c8815331aaa0c4bf43eed5400f116321c4710bd0abc0da30272ef;
// music[257] = 256'ha7ea79f3e8f6cff661031c108d0cae044b08920d300498f7c4f3ebf192ed81f0;
// music[258] = 256'h0b062e1a2d1a8c1679169a109900b2f280f9690b9014b912ab118d16d30eb4f9;
// music[259] = 256'h9cee5fee38ecbde7abf12a0db118330a1bf93ff31f02d915dd17440d6afa04f4;
// music[260] = 256'h8202ce0c3d13730fc5fecf02ca170126662c6d235d10080dfe1d5631bf32a21c;
// music[261] = 256'h8d0b430f1e13e5106412061f3c2e3f2c221e1c12db12bd22392d0c24400e3cf7;
// music[262] = 256'haee8bceafaf496f322ed38eb71e549e174e6d1eb70ebf6e574de8edb5edbc6db;
// music[263] = 256'h62e1e5e6ffe962ea7de743e6e4e4e7e614e9cde664ece9f69a008100e3f3d9ef;
// music[264] = 256'h7ceae6da86cf4fcb3cd209d69fd2bdd0b3ca7cd70eeef3eb7ae581e6bde8d2ea;
// music[265] = 256'h23e6e1e288e510ea13eb84e5dedf05ddb8deb0dd11d929d859d6e2d582d3c1d2;
// music[266] = 256'hadd929db20e05fe079cea1c084ba5db5d4b08fbbaed421da3ade41f06ff5c0f2;
// music[267] = 256'h3cf23bf18aea07dd18d83fe6acf5ccefdae92af2f8f747fc6efc74f9c6f9eff9;
// music[268] = 256'h20fc8bfed1027e04cdfe77fbd8f0a6e202e5adea26eaf7eb2ce313cc09c0dec9;
// music[269] = 256'he4dfa5ecdedc0ec094b490c50bdf5be894e02fd67ed764d873cfb8cb1cc7b8ba;
// music[270] = 256'hebb5ddc832e5d5ea15e628e8eae73ce9dbe774e1eae10de7deeaa8e87fe410ea;
// music[271] = 256'h8ef081f166efeae7d0e617e634d821d332d847d627d023cb3fce94d31fd5e5d5;
// music[272] = 256'h03d353dab2eb2af2a3eaecd8f5ce1fdbc7f02efc56ee68d653cf09de78f45bfa;
// music[273] = 256'h88f8eefb3cf87cfd360e09148b17db1dba1a6710f40986082c0eeb1a2a1a4d06;
// music[274] = 256'h51ef7ceb330098101916b41b421e0d19a30d130f1b0fc901a6fc0aedd5d6d7d5;
// music[275] = 256'h2bdae6df14e77de72fe537e2cde1ffdb4ad291e209fffe0271fb63f48cef67f5;
// music[276] = 256'h91fb3effe0ff0300d3019ef8bef0e9ecc4e114daa9d67bd273cf07dc4ff4d8fc;
// music[277] = 256'hd2f68aef36f1c4f187e085d0d4d451e642ef6af1e7f7f5f76df697f526f18eeb;
// music[278] = 256'h37eb1af392ed0bdb66d2b6da1fec4cf59df94af8bbef90e8abe522eb4aed7cee;
// music[279] = 256'he6f070e34ad980df1bef53fa39edf0d61fcf80d702f25c0ed50dbafc1cf64ef3;
// music[280] = 256'hc6ec6de4c0f0c80b4014d7134611d60b2b09360c19149f05b5f0fcedecf1cef5;
// music[281] = 256'h9df712073f170113ad063afadaf7fef204f63401e7f17be5f2e0bbd387d45ddb;
// music[282] = 256'hc1de13dd6bd97dd962d73ed781d834d963e2b5f85d06f4fa90e649d94ee24ef2;
// music[283] = 256'ha2f453f649f721f6ebe9afd516d6aee77df956fc5ceda0de59dc6deb8efa89fa;
// music[284] = 256'h32f71ff9eff61decb4e13ae325f5ec019400080036fc89f8d8f7c5f9ccfc68fc;
// music[285] = 256'hee0066f719df68d828dd3ae18ee105e2aae327e577f018feb7ffcfed63dbc2de;
// music[286] = 256'h47e2fee880fa3802fd0441081504c4fac1fa710f24257a20720935fffe081e12;
// music[287] = 256'h8c0cc8098c16c51e1f20e122bc20891f8f23cb2a9c24a9018de612ef0302d10d;
// music[288] = 256'h1b116212cc116d0038ed0eea20ed52ee98ed8afbd10bc60a190d4311e90fb90d;
// music[289] = 256'hb50c670c54f909e819ebf5ec4cec33ee33f82efe5ff6abefb4e981f0beff6404;
// music[290] = 256'h9d0498034008be04b6eebfe229e78ee972e42ee936fcb007deffa1eaabdfc3ea;
// music[291] = 256'h57ff1908e1f86ae663e38bef46ff6b032703030392ff05f65aea2aeb87f216fa;
// music[292] = 256'h45f97ee47cda85e3e5e592e42ddf04dae2e7d000e214de1a6411720149f7cfff;
// music[293] = 256'hcf0fa616ca13d80adf082d0799fb88f22bf0caf217f61efc25025c00b1ff26f7;
// music[294] = 256'h06f1ddfd87023cfb79f01de767e8cde9ceec31efacecc3e9f4ea9ffd350ea70b;
// music[295] = 256'hb60773071d05acfb35fab600acfd42fdf1fead0157052605360d000fa40b190e;
// music[296] = 256'h260e521b3928792afa29dd20c020d125d929932a481298fb9af9b2fb41f92ff8;
// music[297] = 256'hef065a10160864024c047c0308f7bff065fade07290c2ffdedf07bf14afbc00d;
// music[298] = 256'h9d1478163a1f73235d209a192217dc111c035ffd9f0dc425cd34ce37f3365d3f;
// music[299] = 256'h0e47ee46914a5f41822c5327c4367d4c8452f642c4310e356248df59d7593a43;
// music[300] = 256'heb373d3d1d3fa33f1a3cb8385b323c323838f028b627bb3a463ed33c293ff343;
// music[301] = 256'h593863236f2345290f298524a92abd3af23ab4386f3cfd3c4a2ec5165115e216;
// music[302] = 256'h62111a1481152c1cb51f3417200fee0ca81422150c16aa29f130582af02a442f;
// music[303] = 256'h9d3126302f33572ba81138065c0ee81f082c1c24a4147109630f6c21b627051d;
// music[304] = 256'hf40abb059e103a1f48252519e70a7208d812901de41c692151275524ad20531d;
// music[305] = 256'h611ced1be01c331a200753fba912ee33223f603eaf3aad35a62cff19e1134e16;
// music[306] = 256'ha7119e14ec16e513c4124012e3122d134e17331d18201c21491bc5112f11a712;
// music[307] = 256'h5803a8f94dfc5dfde410f6221b2195205f20ec221b24df23671d7e0639f9c2f8;
// music[308] = 256'he6f8b8fb5106e11e602730163d016bf60205741af51f1e1c34140f11c519fc21;
// music[309] = 256'hda1fef1fd41f561a0d207628a826ca1f54187617e11aa31ef81d990f1500a504;
// music[310] = 256'he2189a242121aa1d3f21b81f590f6dfe27fcca085b1c3120ae109f0583ff1bf7;
// music[311] = 256'hf3f330f77cfde8fd9403b7198423ec24162bfd25542030197218162d3e371b34;
// music[312] = 256'h0e375c3c583e2739fc35992f631c9a0c4f0e1c16ac1332152a236c2e372d941f;
// music[313] = 256'h4e19a2181511860cd10d5a13de0935f9a1049113d115f1191a19bc0cb8f3efe4;
// music[314] = 256'h00f3da069c0a8d046c042306e60465060909330cb5093403b2fdcbf943fb7bef;
// music[315] = 256'h4ada58d864e51ff746f99be19ecc01ca90cf19ccf9ca14de6beb08e810e3f3de;
// music[316] = 256'h6cd691c4ebba96c3d6d2dedc27cfffb844b640bceebc7cb694bb3dcd20ce89ca;
// music[317] = 256'h3dce98ce1dd0fecd6dcc4fcf27d1dcd00bbf0cada8afdbb07cad52ac46aea1b0;
// music[318] = 256'hfab315c70fd40ecdb6c70ec1d9c3efd9ece9c9e5a8d2b2c539c887c9a2c5bcc5;
// music[319] = 256'hd0cd55d52ddd0eef8ff82eeb74d638d013e107f5c1f5c9eeeeef6beaccdf7de5;
// music[320] = 256'h28e7c5d209ba11b8c3d3e1e661e5f9e378e4a0e4cdd52cc4aec4ecc635ca34cd;
// music[321] = 256'h1cca9ec596c284c593c35bcad8e309f0ffec23eb47eff3e818d386cb51ce7bd0;
// music[322] = 256'hc9d311d3f7d356d174d76ce71ee985e9e1f2bcf908eea0d41ecc5acf46d27cd9;
// music[323] = 256'hcee633f4eeeeb2e038d718d7bce976f612f537f7e0f809fa0dfb4cfb53f5cde1;
// music[324] = 256'h02d78de233f76503abf8efe3f0d81fe12ef72efefaffa312d8184e087bf54df1;
// music[325] = 256'hd3000c0f710ff4013af2bff6c408b918fb17070492f457f260f86dfee7ff49ff;
// music[326] = 256'hf4f866f80e05c1132415d50ab30975fe7ce0b8d471d825dd33e212e293e03be0;
// music[327] = 256'hebe30de5f4e0cfe942fe9c061af5cfddcbd7bbd8d9db20e120e383e568e22eda;
// music[328] = 256'h95d702da58de79debae0c8f16201f60141ffb2fee0f60fe4a7d68fdd51f15ffd;
// music[329] = 256'he9f4f2e37cdd8be7e1f7a3fe0aff8fff75fc3ff672f20ff1b6e733dcd3dc61e0;
// music[330] = 256'h60dc2dd7c4e1a0f55cfa5af63bf6dff823fca1fe1702cd005cfec3fb7feeb6e0;
// music[331] = 256'h73dce4ece20fac16eafda0f325f737f626f472f212f60dfaf3f5b6f211f195fb;
// music[332] = 256'h1417bf23191f741fe121a317100309fba8046318e0244710dbee6be4a6f0e600;
// music[333] = 256'hb707d1090f0ef7121e141d13a60a2ef455e5c7e5d9e6abe78aeab7ed3fe79fe5;
// music[334] = 256'h93f859050305a5062c0980099c09790c4403a9eda2e7def44704a209eefc69ed;
// music[335] = 256'h08ee52ef6eea11eabbe601e42be771eb2ceca3e943f93f10ad11090a6706b502;
// music[336] = 256'hd7f281dfb1e264f6c40531067c039506e70054f1e5e227e746fd59099f08d907;
// music[337] = 256'hfc0aa50413f003e7b4e802e772e4e5e16ee964f9f40c5921ea22481af7163413;
// music[338] = 256'hca113a149318fe0e6af684f0a1feef0f3015d105fcfa31fcf1fb33f674f42104;
// music[339] = 256'he0145714d0ff2cec2cee17ebe4dd8edd18eda0fe32fb5eebace2ffe78efa4f06;
// music[340] = 256'h7f09cb0b550a6cfefce603da7ae589fa7f019efc3501fa047ef8ace580dcebdb;
// music[341] = 256'h0edd35e217e56ae180e0c8edc80086003ef079df52dc8ce11ddf38e7dbfc930a;
// music[342] = 256'h0200c5e304dcbce3ade4a9df10d71bd6d5d8b7e3fbfc7109f7fa50e2e6da0ae1;
// music[343] = 256'h2de140e150eb5bff220831fbc9e74edc08e7c0fb5a06ba07f90413fc91e5a7df;
// music[344] = 256'ha0f700046afdd2f533fd1a140419d10c8e068e0292fc68f9e204271a6c21171c;
// music[345] = 256'h1c19da16c70bacfc43fbcdff25f8d5f53a04e90c630591f2b0e4d1ebf2efd2e5;
// music[346] = 256'h10e635eb5ce91fe98ef25c027405d3f98bef11f2e0069c1da21e290af2f9aafd;
// music[347] = 256'hb805e1042907521aec2c7b2a701260f6aafbd815df1e861b4911cb0dc31a0f2a;
// music[348] = 256'h6b2cb5179801fcfb21fd67fbacf60901a50f0f0ec206db056b0abbffe5ecece9;
// music[349] = 256'h6eeab1eb39ee8feb6cea38f097f8e5f851fb0a0d5c1d201af807aafff9050e0a;
// music[350] = 256'hcf0bea0d9a0dbf0e3f0f0f0e7d18142aca2df629c62c5f30ff325341cb545d55;
// music[351] = 256'h264405355a36bf47d957bf571b47e634dd34794a875c275dcc5cf75c8c5de55e;
// music[352] = 256'hb652cb3eec2c8723c627792bc9262e287e3706410a412b447043734172422746;
// music[353] = 256'h754ae346d746fd481b49014c923af11f2f1dcc21dd215b234023fd24ab247320;
// music[354] = 256'h9d1f572012261827f52334304c3a433a543b053bbb34741fcd10f517242bf941;
// music[355] = 256'h3c42c82e8c1dff1b6e2f353bd83c623f5e3d2939b9343b38b43cda3c143f9933;
// music[356] = 256'h651e03167a21a3308d34a43354311031b7312030463275326e34523d373a3c26;
// music[357] = 256'h951f3a311f45e048c134cf223d22181dda1b2b24362dc72fa725191de116751f;
// music[358] = 256'h52383340ec3eb53d943a673f63430239791cc405b801b80158ff34ffe0143c2e;
// music[359] = 256'h332d10256c212522df227424d925481598054c042a0106ff1b017c065c079609;
// music[360] = 256'hf2184b209919a4179c1ec822f020911e47136105f7ff2e022e0e6214a4146b1a;
// music[361] = 256'h2019440ad4f388ebbbfd8f14641a5305a6e8a0e494f942104114c50c9f0b7f0c;
// music[362] = 256'h200464f692f38dfe2609660a840a240e4e0702f5b4e7d4ed4402490be30a8311;
// music[363] = 256'hb71789123d0067f4c7fd03054a00e2081c23bb312424c70c53024a0027fed0ff;
// music[364] = 256'h8702fb05260acc083a02d2fddb0a65222226c314ec0299fe29060106a7f864fa;
// music[365] = 256'h5b0bd808def99bee0ce6f1e61de54ee698f63c010dfb6ae627d74cdf0bf3b6ff;
// music[366] = 256'hcaf832edcbeba1efe1eeede4b0e817f9d1fef5fd81f921f6a5f535f85df908e6;
// music[367] = 256'hdfd0a1cfc4d4f3d55ed5a4e04eefb2e7abd0e0c2dbc67bcba2c56cc3e8cf00df;
// music[368] = 256'h9ad906c665bed8be23bcafbbb8bd99c084c180bccab688b17db705ccced365ca;
// music[369] = 256'h3cbe05b9e5c3a2cf46d112d1ead2a7d2f5c5e6b055af7fd093f25df39ddfb4cc;
// music[370] = 256'h57ca8ecf7dcc2dd466eb94fcb3f71ee0f7cb46c6f0cb90d122d93ce8cded0eec;
// music[371] = 256'h2eef38f246f1a0f143f3f9df46c576c3cbc637c4ffc2ccc0cfc196c62bd6a8ea;
// music[372] = 256'h1ee978d476c5e5c519ca9bc8a5caa1d020d0e7d2d1e287ee24e801d8f4cb02cb;
// music[373] = 256'h0cced9cf86d823e87feebee427d5e3c9e1ce78e239effcf136f317f303ebfbd6;
// music[374] = 256'hedccecd9a7e9eef0f9f30af7baf443e3f8d18ad2c7d7c3d4acd3dfe052f206f6;
// music[375] = 256'h40f493f8bcf607e7c3d8f9d9a8dba0d227d3cae74bfe6afca6e672d992d6dcd5;
// music[376] = 256'h9ad581db6ceff4fc31022d10ae150a092afab5f6e3fb0df823efc6f7ab0f9c1a;
// music[377] = 256'h600d40f8d6efa4fddd1136168107d1f448f2770046140116dff87ee469ecfbfc;
// music[378] = 256'hbd0c430acbf701ee17eedbec23e731ec9dfd040852091f08a50b840807f581ed;
// music[379] = 256'h3cf3d1f185f056f7d8041109c9fa73ed80ec0fed39e993e7b3e7c6e840edeaee;
// music[380] = 256'hf3ecefe88be678e7bbe796eb7df093f2b8f2a3edfee9d6e654e195e747fb9a08;
// music[381] = 256'hb301b9ecdededae9ac01ce0da6069df366eb7cf3d3fee00462f91ce7afe21be8;
// music[382] = 256'h9feb7dea62f2db0043052e07cd0b3008a906df175724611d80189318ae177217;
// music[383] = 256'h071a721d5a1c581b1c197a1bca1ced0a67ff13ffb6f4d9ee6cf10af6d9fb2cfb;
// music[384] = 256'h5cf588f0e2e91ce0a6dde3e2f4e28ddf0ae685f6c5fc68f256e3d3dbeae7a0fa;
// music[385] = 256'h3801ee037f03e4fccbfcf500effe31fcbcfb45fd31fe4efd5bfe94fd1e00d4ff;
// music[386] = 256'h65edbade31e25af0acff3905ed066305a9fc63f320f1e4f94c04f408e000b2f3;
// music[387] = 256'h97f192eb34e337e552e5afe1acdf64e4bae83de523eb74f452f425f9b6ff99fe;
// music[388] = 256'h58fc4bfc4900360251fea3fbe2fabaffc8fc82e7dedd3be305e675e65ee86ffb;
// music[389] = 256'h1c139a164213a714c317b31749171c1ad61a8318c80ca7fb52f6f1fee810b91e;
// music[390] = 256'hf8220b245a1afa051ef615f9290bd1148212a408bcfadcf9b2fdaffe1d059c05;
// music[391] = 256'hea05a505b2f4d9e393e249f38307f805edf23ae0f2e589fe1d07cb03e202ac02;
// music[392] = 256'h35034006530d26072cef31dfcade2ee1f8e606f6890320fe69eab5df1be4b7ea;
// music[393] = 256'hd5e803e3e9ede3fd9bfd22fa20fad1fc02001f02edff79edb6e045e107de27e1;
// music[394] = 256'h9ae68de838e6bddc99d9e1d81ee12df8d902c1016003d90331fae1e488db2ce8;
// music[395] = 256'hfef8d30146f89be5bcdf51dffee1f2f18d05a516eb1bc2094ff63af9b80a0118;
// music[396] = 256'hc2186e18581fb41c1b0864f5e2f87b0f341e6a1b0015900d6209ea0b76112e0f;
// music[397] = 256'h99f31cd932e095f365fe8cfe5cf19be2ecdec1dda9dd72e402e6fee416ed84fc;
// music[398] = 256'ha409050534fa7cf83ef671f507f97dfc42fd7dff0410f42105206314bf05a3f6;
// music[399] = 256'h54f4f2f7c502011fcd2f582aac26c82726205c0dab00d4fde6f78df3adf440f2;
// music[400] = 256'hd1ea90f11b07100f0d0a9809a509150132f66bf5a2f7fff22ef22805811c801e;
// music[401] = 256'h8919771eec238c1e88122f0eaf0ac005010f642405360a33731d3515982bd547;
// music[402] = 256'h795311507941b637a840f1521d5c34580c59b55ce451693ec4357344425db769;
// music[403] = 256'hd2602c4d94446f4d905d2261e0506936b127163aba4fe049f4342324262b1040;
// music[404] = 256'h474e064eb03d8c3306348d3334336b2d2b29072d2f30d731c031ae2c46267723;
// music[405] = 256'h802d8143c14c853e262d312b33307d2cfb282f2a442b722a48242a21dd21ff21;
// music[406] = 256'hbe233224d1235e1f791c101d411c0c1e3a1a8c127413cf19c8191b17be24a82e;
// music[407] = 256'hbf2d17328830aa2cb1293529752acf24e527d4253b16f00b4205f4014301ff0d;
// music[408] = 256'h3621be2344230d25e22d213c7b3a28345736a43947399a373b38353c423f733c;
// music[409] = 256'h043b6438b2325e313e329737143474224d1502178425592bf02b7a32ac2a251c;
// music[410] = 256'h7b18c41ca4186706f3fb93018f0f5e17a10fe00209fdf00a881b4f190d145612;
// music[411] = 256'h3b10bd123919fd1db61c1d174e1252124e157b18fb175016011735136c11bf0e;
// music[412] = 256'h56ffdef428f68ef71df6f1fb200d03142a0d6a0aa10eec0b3cfb83f36ef7b7f5;
// music[413] = 256'h5cf5fff7c0faeff992f325f0b5f2ea03ee1731192e15d6101b0b5d0bc50daa0f;
// music[414] = 256'h770cfc07ba085f0bf60ef10d440b5e0dd20d040343f4a901ce20312adb1ee90d;
// music[415] = 256'hbc0739122323712f2d28a815ef09620c3c17481b981faa294f2d8d26781d2b18;
// music[416] = 256'hb90f42079b052e10a31d3914f208c60a1207d808c70cdd05b5ffbeff4cfee3f9;
// music[417] = 256'he200910505f315e1f2db4fd9fedcb3e265e123e097e175e19fe13be036dd20db;
// music[418] = 256'h7add75e196de6ee0bbeb68f4f3f90afc39f7f4e5efd1b2cbe5cd25cd47ca4ad3;
// music[419] = 256'h00decadb7fdfe2e4b7e3fde1f8dee4dcc5d5c5d168d161c4a6b813ba49c61dd1;
// music[420] = 256'h56d482d757d4d2ce99cc6eccb9ce75cce1cba8cbb6cacacec0c89fb81baf64b8;
// music[421] = 256'h06cbb6d08bd0add0f6cd06d584e383e4c5d456c67cc7cbd929eabaec98ec19eb;
// music[422] = 256'hc6e50ce1bfe6a2ecdddb5fccadcb26cde9d05ad505e8cdf7cae994dc5bdbc7d7;
// music[423] = 256'h4fd4b9d6e4da29dba5dd45d744c828c7aaca5ccac8c96ec8becc79d155d120d1;
// music[424] = 256'hced1ddd60adddddd3cdc02d4cecf35e347f886fb2af73cf3ffefa9e32ed946de;
// music[425] = 256'hb1e77df08df01ee7bfe0fae458f202f5ddf07cf3d9f54cf725f74af8ccf41ee6;
// music[426] = 256'hc7e09eec4ffc3efefbf703fb89ff55020103dbfed0fdaffd5bfd65fdc6febaff;
// music[427] = 256'h6df34ae3c9e42bf4d7021602fbf1e7e7ebea57f559ff18fd3dfdbd02d100b7ff;
// music[428] = 256'h8efa94fcf5104c1d1220e421dd21b4193e075e004e0201fe1ffb43059918981c;
// music[429] = 256'h6a15bb17b21af81071032c03830480ff34fad4eb73ddc7da25ddd2de16df91e1;
// music[430] = 256'h51e02ae264f123fd5bfd52fca7fe12ff06fd29ff37fa6de7fedc7ee71ff785fc;
// music[431] = 256'h7ff465e76ee016e4ebf170f8cded64e134dc36e80efcde003cff07fdbaf9a6fa;
// music[432] = 256'h1ffb0ef883eca6de9edf9defbffec4ff77fa7dfaa7f92ded34dc9fdcc6ec75f8;
// music[433] = 256'h12fa07f95ff912f271e146d89ed939d873d6a8d922dd4ddfb5def4e042e19fdb;
// music[434] = 256'hbce43df100f311f5fdf4c6fd6b0cb80d350d98132616b20645f3eff18ef5d1f1;
// music[435] = 256'h90f10a017513f510c6fc35ec8aeb3cee4ef129f64bf59af86ff65be5e9d9d8dc;
// music[436] = 256'h87ea81f3bff65dfa4ef6a4f185f2f0f75dfb6df989fa90f904fb6bfc6fee66dd;
// music[437] = 256'hb9d9f3e6bdf6fbf9edf089e38ce31cee5ef5bef3a7e6e1dd2fdf9fdee4d757d7;
// music[438] = 256'hc2e7cff996fa28ebbede72dcc1d9d6d873da0fdecddeffe326f8b901c6ff85fe;
// music[439] = 256'h98f76df488f26bf53cfbeafbc4fef7f2f6e066dfdbe08ce248e4c2e10edc9cd9;
// music[440] = 256'heddd5fe224e625e4e8dd47dbe8e766073f130e0465fb0ffe93fe76f4fdf39b05;
// music[441] = 256'h6910500fc210841ad91a880888f8e8fa830afc13c714f2145016ac166115d11a;
// music[442] = 256'h0011f8ece4dc61ecc6fc91fed1f876f742faa9fdbeff96ff7ffd86fe91fe7cf0;
// music[443] = 256'hf5e6c9ec18ee97e587e2faf390074304a7f293e558eba2fc6306e7fec8eaa5df;
// music[444] = 256'hf1e1aae230e124e862f6a7fefb00c106650989faa0e7a5e637eb07e6dedfdbe9;
// music[445] = 256'hedfd8605ec05cd07d0069d0251fe5efe8ff692ea3febf8f2ccffec0262f35be9;
// music[446] = 256'h55e70fe4eae1b4e292e452e4cae6cbe9c2e8a8ed60fe8b0d4a04cdf145f9df0e;
// music[447] = 256'hc11e4027131e6309b8015911ec269f2b69216d1464131623902f7d2d8a224a1d;
// music[448] = 256'hdf1e40171710700fdd0655fb6df96dfb68f1c3ee9b007505a5008f07a60c9c08;
// music[449] = 256'h100847112d0cd9f5e3e9c7e950f138f927fba9ff0502a601a0040307fd074b08;
// music[450] = 256'hb608430bd60dae0c99101e19a3140b11d41eab2367120e07b112ae287c39d435;
// music[451] = 256'h71277127772746164902bcfec10e701c9a1a9a13d10f1d0955fba4f17df62506;
// music[452] = 256'h010e4a0d7b1356174319d81d8518850fdc0c2e0f44122d16be1bc41837155817;
// music[453] = 256'hd90de70107047206db098b199424ff24f02b963cf5496a4525365e2da72c432d;
// music[454] = 256'he42b0b334246d553074da63b8034e435c933602f263c3b56535b4c56054d7e35;
// music[455] = 256'h012e5e35f73c284733470c3fae366e368b3b65348a248d1e66290036aa3bad40;
// music[456] = 256'hbb454e430a2e6a1c5a1ebb1e7f181d191e2d5941403b28285219fe16c5193c1a;
// music[457] = 256'h18227632873b402e651b1f15cb1dab307e34c4306f32c72f6a2fac2f0830082f;
// music[458] = 256'h102d0f2dc51e6e0fc80e4f119f106910661f6e2e9b28e7140103b30632183224;
// music[459] = 256'h20219d11ec0a090bd90687ff9a03d418fb251c1f970a7602c314ac1f741f861f;
// music[460] = 256'h0f1a941770212a33eb37e031c230d02e4c303635343500285d129a0fd61e2930;
// music[461] = 256'h6034912401179412d912090ee9fdf4f766f997fdc2064a031e0234104216850c;
// music[462] = 256'ha1ffe4fd670560064bfdbcfcb70e6b1c891b5019cc1439081ef8b4f47703b311;
// music[463] = 256'h5918651b4a1d021c4909edf354f340f9a5f926f7ebf78df9b0f9950821166b10;
// music[464] = 256'h420bda0a010cd30d4c0e760a11fd19f880fd87fcbbf79ef81c07a8147c121605;
// music[465] = 256'hc6f611fb0e0b4d11470a35fcecf46bf3a8f13ef3f900aa15f117fe0822f7d6f0;
// music[466] = 256'h6c01f10e9f167c27942fc2260b14b005140dc12092282621471cee1f97205e14;
// music[467] = 256'h2d074c0aca165b22a61e2f0bed02690442052f064f047105b7ff15f51ef4e5f1;
// music[468] = 256'h6df6200a17161d091ef041e98cece5e99eeb6aecbee83ce7a0f13a04e00256f2;
// music[469] = 256'h14e9fae894e941e47be8f5f73a0396ffefeb11e319ebacee46eb41ea51eddeea;
// music[470] = 256'h3def93fba8f98ef14aefd1f438f83df3c7f126e50ed1b7cdfbd1a9d184cd6ad3;
// music[471] = 256'h58e0a9e18dde26e00ee202d948caf8c5dec255bf21c5b9d2badec0d93fc824be;
// music[472] = 256'he4bfe0c2fcbe18c052cfe9d9e8d723d940db80daf8d77ed1c3d9ddec21f217ee;
// music[473] = 256'h8de91fe909e528d80bd70de5a3f228f4dce428d3c8d03cde47ed55f051e58fd8;
// music[474] = 256'hfbd5ebe1b6f651f35bd4c2c3fcc3f1c272c044c37ad420e432e172d2fec6a3cd;
// music[475] = 256'hf1dd75e7fae1c0d1c0ceabd344cdb3c714cc47d789dfb0d976cff9ccbfcc25c9;
// music[476] = 256'h45c8faca2acc27ce3cd152d4f6d654d695d0c9c8dec8f8cea4d21bd3ebcd29cd;
// music[477] = 256'h18dc38ee09ef2edecad268d3a0d499d404d24bd1c1d549da04dd83daa4db30e9;
// music[478] = 256'h1df208eaa8da1cd5ecda52dd8ddd7fe6d4f21cf633f51cf88cf72ff992fcabf6;
// music[479] = 256'h6bf92707c40cb90c2f0e820e040aa30b320f3c0329f6d3f2a1f277f003f21802;
// music[480] = 256'h800dd60de90dab0bf30c640f7611d30a22f822f494f1fde341e190e993f95d00;
// music[481] = 256'h10f3ebe40edf40e8adf903025a040f04240051fa3bf702fb74ff38ffccfce5fa;
// music[482] = 256'h0efcb8fb18ef4ce001e4a2f4230145fff2eef8e0dde4cef4e5fe7bfee8fd6000;
// music[483] = 256'h01fc6dec0ee241e873f53cfdacf5a6e7f2e329e4fce1b4df73de0addf8dab1e8;
// music[484] = 256'h58ffbb041b03a10094f834f59ef7c4fb3bfb49f8bdf436e6eddb17df5be17ae1;
// music[485] = 256'h0de04be04fe29ce12be31be218e4cbfbb713c60c1efae9f6dcfa7cfb70fa03f8;
// music[486] = 256'he6f4bff349fdcf0d4011500c970d450eaf07bafac3f5b602530fbe11940efe0d;
// music[487] = 256'h77104e0617fc78fa36ed8cddbadef7ebf7f55ff9c4fd54000bfecdf7e0f53ff5;
// music[488] = 256'h4beb4de509e632e4fbdf55e4fcf7cffe0ff8eef9fefdf3f90de9b1df6ae9d4f4;
// music[489] = 256'he6fa36f274e486dfb2debcdfa2e12ced65faa7fc70fd34fe3dfae9e96adc36e2;
// music[490] = 256'h3be675e3e4e8fcf96c0546fe6af7fdf837f699e883dd9fe584f61a01ddfb2de9;
// music[491] = 256'hbedf11eab4fb1304eef8d3e338de12e671e837e880e595e2b2e35beb0c037514;
// music[492] = 256'h9f0b06fdfbf90f06b2138b118e04c0fcbd05c61a9325311d190d17016806ee19;
// music[493] = 256'h23269b22801072033506a2070709cc07cdf88dec4fef5bf747fa02fa21f574ee;
// music[494] = 256'ha7f75e09bd0c780531060e0dbf0543f7c5f242f2e5f4a1f90ff947faf7fee7fe;
// music[495] = 256'h62f934f318f133f20ef474f49af10cf08cf111f345f4c1f4d1ef9aef00fe2f06;
// music[496] = 256'h9f06dd0a850956097509b8066f0842081407e8ff4cf301f2d5faf404290343f6;
// music[497] = 256'he6e999e84bfb980ddb0f900b85071d06290477046f07ca08d806be0296fea1fc;
// music[498] = 256'h2302be06ce0a150ecc05d70a1713ad010af417fd9d0d2d0f2009f30d890f7e0e;
// music[499] = 256'h9c14d61e271f730feb0229f982f30cf7daf8bbf9b1f645f484f40df498004908;
// music[500] = 256'h090014fdb3fa51f5f7f84e03d109fd07a805870464ffebfbd6fa83fd23080807;
// music[501] = 256'h13f583eaf9eed1f799fbbe03a1183e25b0210c1d6119a2104f0677054a0bd30b;
// music[502] = 256'h7b0f5b19b61e4d2457275a24a521b61540076208ce1262159d0cb90679057805;
// music[503] = 256'hc5070c07610786070207f106e106e20cd908e8f653eb95ec32fc9d0b1b0d4503;
// music[504] = 256'h4afbbc01b30c42132012e808e1037502cefed9ff500c391c202c5639693dc43e;
// music[505] = 256'h2f379b2bac2e9032d32ea32d7f3bdf4b6b4ae948984c9e4c894ba249c548a745;
// music[506] = 256'h8e49004e2e43813c063da5351728ab217c249a238a24772697225621031fd31e;
// music[507] = 256'h6c2a8e39b23d71300320261f142a63354d3a992d481984177c26e135ed343121;
// music[508] = 256'h6210801238255b333a32d9315f35aa33dd2eb42b75231d14ed0a18139525f32f;
// music[509] = 256'h8d3105304e2bf02a552a0e260c2361258c2bd121770c3d0126fee801d80aa913;
// music[510] = 256'h9316fc0ea104b3fec200b509530f8a0d1f080dffe9f74bfc8901170856189e1e;
// music[511] = 256'h551938185b1fe5298923b313bd113214cf142c1cfc274e2d422b3b2d9930052c;
// music[512] = 256'h4a285a293b22a313350f801c0a2c7c2c83273427e826312aea299d1bcf0fdb11;
// music[513] = 256'h8418021db91c09182614b012720ec0010ff5bdf8480a6f182e15b10234f6ddfc;
// music[514] = 256'h830df7164d13c706c3fad1ff4a0f7c1551173219db16bf0b4afb3cf607f91ff6;
// music[515] = 256'h7bf50201fc0fb7132511c30eef0851097613dd179b167f1da524f521a21f2f1b;
// music[516] = 256'h580ebc05d905cf070508890554044a069b065f07f70a300be8065800fefc5fff;
// music[517] = 256'hbc007207ca15611b6913e30758053211701f4e244c256321be1855201b2ec42f;
// music[518] = 256'hb53483389b33e731f8310732db32bb31f02aa11bdb0e6114dd26e0318032a531;
// music[519] = 256'ha72eab2c8c2fa82e9c229e16d513f60ff60ce114b516ef064df818f36aef93ed;
// music[520] = 256'h40ef18f4bcf5d6ef2ce9b6e632eb11f052f3cafeb908d308a4062e08150a0606;
// music[521] = 256'h1c04e30079f46ee6d1d9cfd4d3d1aed222e4edebade359e07cdd6edcf2dce0d7;
// music[522] = 256'h9dd35bd3a7d5c5d295c490baffc22dcf44ce99c90acd26d359d219cccfc6a7c3;
// music[523] = 256'hd7c779ce05c8b5b971b200b9b9c306c407c3a4c706c8f4bd19aeefab0fbaa1c4;
// music[524] = 256'h4ec71fc623c235c70bd83fdf53d8a7d482d6cfd96fde12e4fee0b4d044c991cc;
// music[525] = 256'h77ca12cbbdd473e0e3e102dc14e0e2e5d1e4cee653e35fce51bbceba01bf8fbf;
// music[526] = 256'h54c19dc71cd173d1b1c7c1c01abf32bff8bf04c3bec6b5c5c6c233c17ebfb9c7;
// music[527] = 256'hc5dc16e9b6e42fde14dbb5d561cff0cc3cd065d978dbcfd1f4c775c40dd2c9e2;
// music[528] = 256'ha0e15edf59e449e7e6dd8ac9b6c35bd085dc16dec2d586cebad227d7f3cf53cf;
// music[529] = 256'h27db61e324e626e6fae8dee9b8e59de43bdf59d4a6cf48d7fde637f13bec51da;
// music[530] = 256'hd2d079d2fed1bad154d15ad24cd40fdceaecb2f148f264fe220576fcfeef72ec;
// music[531] = 256'hb9eaf7e842ee76f4e3f5a0f159f547045409c1fd01ee38ec2bfacc081e0b5706;
// music[532] = 256'h5609a50165e90adeb9df25e15fe089e0e4dffeda91e265f59bfd8afaf4f4aff3;
// music[533] = 256'h4ff481f5c5f650eb24dda7dc72e03adea6daf0e688f9b3fb16f9c8f866f452e7;
// music[534] = 256'h0ad9dbdb5be28fe24be4e0e131df82df55e90afc93fee6f086e3e8e064ebb0f2;
// music[535] = 256'hc1f243f6bbf979f11ee09ed487dbd5f05bfb1bf889f8f8fa91f574e5aedb6ee5;
// music[536] = 256'h6cf424fb19f2a4e30ae298ed05fc93fb45ef6be88de8b5f204fb6ef47cf7ba0d;
// music[537] = 256'ha6134900e5f46bf7bef8aef751f5c6f333f2fdf695071513390e60fe76f5d3f7;
// music[538] = 256'h1ff6b3f520fedc0e971abe0947f738fd4bff3ff44cf3aafa39fa1cf90df830f3;
// music[539] = 256'h3af5c6f813faadf91bf687f645fa5c05f911740ebe0043f736fbd10837135215;
// music[540] = 256'h32140d14c30a18fbd1f287f130f250f6d504ba14771625066aef54ea9af138f6;
// music[541] = 256'h1dfa5c02060b7a0636034b0ade0c370d8408ae031105bb093e0f980b8d0ab708;
// music[542] = 256'hbaf643ed31f122f322f015ed43ed46e9c0ec2e011312990fd5fbc9ea1aeedc00;
// music[543] = 256'h1812460fb0f994e9dce5a3e7deecbdf4a903ae0be40015f309ec3af517039704;
// music[544] = 256'h5e06460aa30b31fd56e29adaacddbbdf44e183dd0bdd8edebfe1bde418e3dfe5;
// music[545] = 256'he0ebe6f0dbf2f0ee2fe92ee64ae83aedabeebbeb36f03ff636f2b3ed78ebf7ed;
// music[546] = 256'h44ef63ea8aeb91e95ae77bedf5f067ef97ed24fb2f0c4c0b55092b04bafa3cfe;
// music[547] = 256'h2209b310920e97048afef000ff08d60b19021cf7a3f5eef843fee3042b0a580c;
// music[548] = 256'hcd0af4055f0035046b073cfd59fbf50069000001ef02ee041f039e02700647fe;
// music[549] = 256'h3ffa6c0619090504aa05860402fd39f7e6f86efd87ffd80698080cf72fe8d7e4;
// music[550] = 256'h1ce5e0e720e42fdbd2d7b9dcd9e5eaea4ce88be646ef91f8e2f945f56def02ef;
// music[551] = 256'h65eaaee323e547e843e7c3db97dab7ed2cf770f681edc1df39e360ed77f0f6f0;
// music[552] = 256'h02f191f1e2ef6ced3ceb3eea9cf147fdc0fc24f440f11bf127fc32117012a308;
// music[553] = 256'h7a0b360d400d2e134414cf190b17c5fe13fa150090fc8106b609e5046003acfb;
// music[554] = 256'h1afdfdf7e7f0eb015707e0013308890819071008d104f5086b13f0154f12c014;
// music[555] = 256'h5b12a107f0112823362298204e18e20f2118581e83249b276e1fd71be71e6329;
// music[556] = 256'hac321e33273539384239ad34342f70293c1fec227130dd37e33ced3be0366238;
// music[557] = 256'h7b3d0237a929e5260f2f5f362d3473354b3a37384f3c4539a929c124bc294031;
// music[558] = 256'h59320d2d4e2ed63053328c369f32ac22631b282289290931b8362737373a7341;
// music[559] = 256'he539e124cf24172fb52bed2957327e3fd447464808446141ed40a93a763d593f;
// music[560] = 256'hd736ee3ba03f564124434539123abb350c2b4731ba32533718433344a242603b;
// music[561] = 256'h18325930ff29501fe21e392d713d2f41cf3a13314e269721b229233af943bf3d;
// music[562] = 256'h9c2fdd2ebb3f2349a244a33d383a1e43ff45513d8f3294199c0f53190d122e0e;
// music[563] = 256'h640f640aca139119d00ef007bcfd5eee98ed89f3acf762027a060cfbc9ec70e5;
// music[564] = 256'he5e5dae90fe7a3e0c1e576e671de73e2f9de50d399d55dd905dc24e602e6b8d4;
// music[565] = 256'hc3cff8d59cd5d1dcd6db8dcc81c713cac7d042d720daf2db30de07e16dd8f5ce;
// music[566] = 256'hb9ca0cc527cc1ad552d261caddc0afbd76c2a2c874ce2ada74e088d722d49cd0;
// music[567] = 256'h9cc9d4d10edb8cddcbdff9dac3d9b2de0bd678c9e1c9becd29ce78c88fc6c7c8;
// music[568] = 256'h5bbf5cbbcfbdadbc3ccbd5d84cd5cdd1c6d01ecfbfcc6bcdd5d414dbacd85fd2;
// music[569] = 256'h3dd22dd4a0d6dbd855d2dad3ade18ae3e0dabed549db5de374dcf7d217d79ddf;
// music[570] = 256'h8ce3bbe57ce515db33d4d1d9cfdb40dba9dac0d7dad9aee079e9fae591d487d0;
// music[571] = 256'h40df55eceae76fe07ae81ceb68df0fd8f2dc45e922ee5dedb1ef18e5d9d63ddd;
// music[572] = 256'h00e564e0c0e0b4e84fef78f7810264048f00a90080ff22037f081c0426002000;
// music[573] = 256'h9802e4027efaf2f763fd62fd8a01560996037200bc0761035ffc43ffbc05cd09;
// music[574] = 256'h8e04e1003508b612ae18bc175712cb07d101e90682093701dcfa1a04470b920a;
// music[575] = 256'h0d0dbd08ff04480a6e0b0f06eb0a1c17240590e8a8e969f0ffefbef271f535f1;
// music[576] = 256'h4fe940e7b5e438e8c7f548f84dec12e575edaaf60ff42eec44e437e4b3eebef8;
// music[577] = 256'h87fc4b027afc13e89ae5c4e81ee89ef0daed44eb0fede7e631e775e3bae1eceb;
// music[578] = 256'hdaf0a7f4c3f49eea0adf1ce1d9f001f7c0fbe7084c0b5105c506130ca60b600b;
// music[579] = 256'he903e7f247f2d6f803feea06ba04f9ffb7f795ead8f0beff3e003ef45cf1f4ff;
// music[580] = 256'h860c270bd2fe29fd4b055a07780d840eb50d9b15f619561fef16e507440dbb15;
// music[581] = 256'h7c1ee524a321e61dc5188c23f1339a2e3829bf2a5e2ac02c1c2eb72e2a296825;
// music[582] = 256'h1733a735012ba233d63d3f3be536ca333936bf34a930c734e3355030942d5a33;
// music[583] = 256'h3538e535ef346535f63602336a2c8a365043d63baa2bd42bc437f03b6f3b9834;
// music[584] = 256'h87321f38fe2a99212c2bf52e3132f633fd2dcc29ca269527b7371f4d664dbd49;
// music[585] = 256'hc851584306372c535566115c1458c75eee6312606857ac529c4dcf510d5de658;
// music[586] = 256'h9450864f4f51ca537b4eb64f6655c44a454ae2548150ef4fab503846234ac950;
// music[587] = 256'h8946df49b35073445848c9524d46f93e183ff43d78466246f43a6533a72dbf30;
// music[588] = 256'he83675350738fd3931387f370b28a913951244190717e60de907a108a40fb712;
// music[589] = 256'hf50477f87ff663faa806f106270189ffeff030e720e8d6e998ea50e309e877e8;
// music[590] = 256'h80d679d788da22d667ddffdf08e0b8d928c480b718bae1bcd4ba81ba91bb11be;
// music[591] = 256'hdec0f7b750b2a8b7cab48baecbab37adf6b1f5b411b7b0b275b158bb41bfbdbd;
// music[592] = 256'h0fbcdbb648b400b73cba6cb838b433b9c7c259c0dcbc99bf55bd8cbf22c061ba;
// music[593] = 256'h63c029c566c3f0c0ebbdcbc193c41dc725c844c8cbd158cfc8c442c40ac7c1cb;
// music[594] = 256'h32ce4bd130d22ecd49ca1ac83fcc3ed3d7dad9df85d8dfd754dc92dcabd835cb;
// music[595] = 256'hf8ca48d4a1d9ece511e86ae0ccdefdd5c6c9e2d384e4a6e12cdc60d739d14ddb;
// music[596] = 256'ha9e6b2e400df94d928d773dcb7e2b6e179df28e2c7e50be43ce2c2e2bfdb62d8;
// music[597] = 256'hb8d924dc0be5fae69dec02f09bde30d8d6df25ebe6f798f5c3f0e1ead4dc0ddb;
// music[598] = 256'h9de849fc4d0d920f890db40f72057ff932febf031d042804d3037a0116027c0a;
// music[599] = 256'h300b67088e0771ff10009b065b06640497049008f9061a04cd083c0c7f0d6a0b;
// music[600] = 256'hb10362ff490a0618b715b20e2e09b0fb28f54e0259087606f8109d0a2a01a70c;
// music[601] = 256'h5a0bcd0b3b128f06ecf78aea0eecf6f6cbf138ed8be91ee3eae8b0ef4bf226f7;
// music[602] = 256'hc3f341ea60eb60ef66ed3fe8adde6ae133f00bf12fea86eaceef40f91e025903;
// music[603] = 256'h01fda0f173e928f000fcd8f85ceb71e3b4e23ce5c4e8abea07eb82ea09ed18ee;
// music[604] = 256'h05e2aedb8ee8fef6d9043a11590f2d0128f822ff6c08930765012e0096020b00;
// music[605] = 256'h4ffa5ef189efc5f78af952fdbdff0bfb1cff4f05c407e1ff5ef4ddfc5505b006;
// music[606] = 256'h000f9610320f68153c184513e7128f1b3120231d421c83226623a61d4827cd33;
// music[607] = 256'hf22f162a6e268f261d2eb235783930370733982fbb33aa48e3579055064f1c4b;
// music[608] = 256'h1152765488471348025266504656fb5e35586957f5524b47385283547348b14b;
// music[609] = 256'hbc4d5053bf568251f656fa53e24d4d520c4f014a654453401e48be4e194c2645;
// music[610] = 256'hb8407b45824bb745993c133c663f17423d47544f774e9b43923b523bf24bbb5d;
// music[611] = 256'h955935540554274dbd4fa3585e5758584259f14fa44520417b4cc052c947864a;
// music[612] = 256'hcd4ccb43c63f0f3e9648ea4fdd47214420423b3fa13c5938e23c974684464c45;
// music[613] = 256'h3247bf3aae3234359d2d522abc293c23cb1f1b1cb81a271a6b1ba91fc920df1f;
// music[614] = 256'h061cad157006a2f539f291ecd2eb92f8fafa55f7a3f2b8e41fe19de212d7bcd7;
// music[615] = 256'ha6e058dce3dcf0df12de3bdecfd6ebcaecc673c7d3c36dbff4c0d6c69ecc27c8;
// music[616] = 256'h36be80ba90bd9cc4a4c06ab702b50eb503bd5cbfa7baf5bdbdb9f9b370b90cbe;
// music[617] = 256'h6db9d8b0d8b613bc06b054ad7eb416bacabdf8b97ab9bdbbceb703b422b4f4b8;
// music[618] = 256'h72baa5b78aba08baf2b391b7d1bd7eb857b4e9b64eb982c0a7c5d1c257c180be;
// music[619] = 256'hc2b721b986c8ded5a5d5a3d01fcb94c03bba32c60bd3a0d232cf18c906cabdce;
// music[620] = 256'h6dcb37cf0ed440d107d3d8d30dcc08cc3fd4b1d2c9d63cdc62d5c4d70ed844d8;
// music[621] = 256'h5fe313e657e209d986d0d3cf62d2a6d993db9bdd4edfade14be2b6d056cab7d4;
// music[622] = 256'h61dd36e85ce6eae2a2e319dd06d951dd6ee28cdd04dcb7df8ee38eef63ec56e2;
// music[623] = 256'hd5e05bdc77df3fe69eeaf3eb9de7f8e37ee06be180df94e68b026a0bd902d102;
// music[624] = 256'h15007ffaf1f8aefbf10079073f0c0a0bdc1010145c01e8f6d5ff6405a608bb09;
// music[625] = 256'h200b890fa90f2b0eb2033bf92bfff406ac0a74073d053d0d7909feff8e01f200;
// music[626] = 256'h20fe54063115ae16030ebc0eb90ee30167fbf9049d0e04107e0dc30b8b0a3504;
// music[627] = 256'he4f766f094f286ecfee613f0b1f0adeeb0ecdce025e4bdec57ecddf0baf4a2f8;
// music[628] = 256'h68fcbff131e23ee6cdf4edf64ef8dbf953f31bf258f195ec92ec4eefeff84b01;
// music[629] = 256'h57fbe8f4a8f078e6fae128ea76f07feac5ead7f478f012e1a9e019ef12f6d5fe;
// music[630] = 256'h100afe030008110d370a32150e0ca700bf044bffbf0ea61cb012bc125f189d16;
// music[631] = 256'h6c11e211f11241190a25c31a8414ee1bfc192a1af415fb105d1b622a3c323631;
// music[632] = 256'he12f582d9d2e2b37f4371239cd3ecc3802329f358038173ea3456446564ab250;
// music[633] = 256'h1b52cb4e134c2b4e484e7d4fcd4b8f46064f6950204da24f7e4a424d9e562551;
// music[634] = 256'h144d8253564f934c9d501b455342ca4bab4e7a53334aae42e048434381434b47;
// music[635] = 256'ha93e253cdf3e68445949db42bd3cdf39cc36bb3b743bca3ac944f543a642c642;
// music[636] = 256'hf0357a34cb3421334d3f82374a230822e219e818c535f03cfe2f0d35fe31c630;
// music[637] = 256'h763d4c3cd23c8a3d3630ce293c2a7c2bd22e912ec22a9627382b5a336733a62b;
// music[638] = 256'h9623bb1d171fcf24a827c72bdf2d30272522a828c02e252e3c2e282bde23081d;
// music[639] = 256'h981b8e1d6017cb146e191d1d0f23bd25a6275521f4130e18b619820564f4a2fb;
// music[640] = 256'h5409260451f984eec9e6dfeb0aeb84e991ee9fe84fe28be1f7df68e036da8fd2;
// music[641] = 256'h71cfbec721c90ad014cb44caa6ced1cc62cac6ca2acbccc6c3beedb84dbd75c2;
// music[642] = 256'hb4bfebc09bba4cb23dbbb8c354c4ffbb2fb384b4dbb515bbc4bf26ba41b455b5;
// music[643] = 256'hdbb7bab578bad1bfc5bc95b906b681b5d9b270b4cac1bac4c7c356c5e1bf82b8;
// music[644] = 256'h71b2c9b465bfadc5d6c224c272c5ddc28ac773cac0c368c40dc355c6e6ca30c4;
// music[645] = 256'h74c751c8d6c521cdadc8ccc564ceb3cf64cedcce5cce89cf0fd39bd450d370d0;
// music[646] = 256'hdccc05d36bd77bcf92d0b7d862dbe6d9ecd27bcd71d37adcaed8a4d845e026db;
// music[647] = 256'h4bdb98dbe9d78de537e806dc0fd9cbdb88de6cdac4de6ce5f4dccede91e530df;
// music[648] = 256'hdddc90db9ad5cfdb92e481e278e4cee4d9e422e9cadfefdab9e5e0eab2e588de;
// music[649] = 256'h2cdcb1d973ddafe652ecb6f094e9a2ea3ffdbe06c8098d087805d0ff60f80500;
// music[650] = 256'h69058603e7030204a90bb80edc084605c004fd093f0ac705ef06d6068e036005;
// music[651] = 256'hee0aa30b6d09e307b207030a2d089106c306aa04ba0b561100093c064d065605;
// music[652] = 256'hce0e1d128710b5143f11a60d970b4408aa0b63123d154902bcec96efeff0b2f0;
// music[653] = 256'h94f6aff915fadbf629f7ccf27fec86ea38ed49089d16f00812085c07b207d50f;
// music[654] = 256'ha10c360ba413f512e3091c0e3013b80d990eda0e5f137716390c96098605b7fd;
// music[655] = 256'ha6002504090709064a06d20c710876fc91fd5006d10a4013d319d31c0622661c;
// music[656] = 256'hd71cfe21a7182a19ca1f721ff51d05123906c20a0414e5128d0e9e0f88103711;
// music[657] = 256'h5c118413e7150b16d51abb1c381967153813071b8124ec2624268c249925842a;
// music[658] = 256'h032e9e2efb3289348432d1389a3b233ade3a3336a532c134753e284bd24b1049;
// music[659] = 256'he645d13aab3aaa445b3d5231262f9728b425592a8c29c12ab0315432162c312a;
// music[660] = 256'h6b298a28102c8026ab21892af02b3e25fe223325b12add2ea52f462b2f275628;
// music[661] = 256'h9a2622281d2fe22cc328ad2980265c229f214025a429362ac32c5d2977238c27;
// music[662] = 256'h6521d018a5205f200a1b5127ac3770396e345b38cf3b9e387a3a6038a2304d34;
// music[663] = 256'h473a4934582c942bd02cb52af5289230bc3a6f387e337430a926cc225a27592a;
// music[664] = 256'h902a41280225e31b9f1a75296d29521fbe20ec1f281fe5248c23031f9e1cc415;
// music[665] = 256'h1d12b012bc15ec1f8e22e01d881a6217c916cd0889f995fbb5f7e9f08eef75eb;
// music[666] = 256'ha8e9e8eae7ed2aeb6de62feaf4e817e00fdc48ddd9dabfd4fdd57ed550cdb3cc;
// music[667] = 256'h3ad1ced015cef9cce8cd64cb6fc73ac7c6c381bee2c0dac716c77fbe42bfcec1;
// music[668] = 256'he7b8c4b79abd40ba91b7f1b9e2b93cb96bb9f9b714b72fb501b4d0b8f4b9a1b4;
// music[669] = 256'hedb5f8ba91b84fb737bc66b941b245b387bd0fc7efc279bb6cbd59c13bbfd9bf;
// music[670] = 256'h04c9d0c6f7c0cac35cc3e8c6b7c849c7d7cbbdca35c7a6c4b9c9f6cf4ac8a4c6;
// music[671] = 256'h98c9cbc941ce8fcf69cf86ca23c62ac9c3cebed613d6bdd3e3d4dad3bbdba6e0;
// music[672] = 256'hd4dde6ddebd927d690d669d644d68ad8d2db4ade7ce18adf5bda50d8fbd28ad1;
// music[673] = 256'h5bdbe0e204dfdcda2de002dfced446d6c4dc1ae208e88ae2b3df96e601e824ea;
// music[674] = 256'h49ea4fe599e3aae600f03def6fe47de4cae764ebe2f1f2f226f010edfbe95ae8;
// music[675] = 256'h63e9e5e613e5c4f43706c2082b09b309ef061604f3069b106f12d30bc108610a;
// music[676] = 256'hd0111b147b0bec095b0e600dcd0aef0ed71d3c28f824e6226b2523263725db23;
// music[677] = 256'h5826002c5028511f7a218026b625112711245a1c3f208625e620a32294254424;
// music[678] = 256'h4727b121fe1d1d26f8241a248022d2101e0694096a0c3f0eb10ce709c10a3d09;
// music[679] = 256'hc10a6710510acc025e0403048507ce0dcc063afa77fb98043408770c1c0ca508;
// music[680] = 256'h870ee9095203500a6a04bd01290bdf0293fb8afe4cfc77fa2af5a4f356fad2fb;
// music[681] = 256'h6202070916fc81eef1f360fd2001330922121c19a81e0d1bbc18341ad416e713;
// music[682] = 256'ha611ea13a1162c07e0ed54e612ee6bed5eee8ef85efbddfccafdabfa61fe2102;
// music[683] = 256'h52ff76fc01002c056305e608780b0806b506040e5f0e450c0b137619e314fd12;
// music[684] = 256'h5d1ad21a60185a1c891e23257629b6235626e128c329692d35258223c729132a;
// music[685] = 256'h8f2f2331e82bb0282a28992b5c2c482ee031cd317832b230aa2c652b942d322c;
// music[686] = 256'hcf259f2908306a2e8a2b45277f28762ea12b4f248524d727ca260428cf27ac26;
// music[687] = 256'h8e2a1f2ab5291926be1f3a21481e1f211e27241e1b1d9a226b20ab1f97220f21;
// music[688] = 256'h101cf72749382e378e31cd2c52317f3830375639a435e92e3730062fb12ec02e;
// music[689] = 256'hcc2e492fdf2bac2f2b31742a902ebe318e2d972f2a2d73261128bd2702231827;
// music[690] = 256'h2c2e302dd32c952b2b21171e4e243820cd18931a4a1cfd18841aaf212a206a1a;
// music[691] = 256'hd01e911fe71a211baf0f61fc77f48cf6a0fbbaf851f5e4f4b3ecc5e771e901ea;
// music[692] = 256'h5ae6cae058e0c0dc18d70ad63dd81dd9c4d449d565d512d2c4d08acd0dd404d6;
// music[693] = 256'hffca32c6d4c15cc233c58ec070c3e1c8d4c44fc2c8c3f7babbb473bbc7bb6abb;
// music[694] = 256'hb6bcc1b92bb79fb61dbd16bdcab974bc13b816ba49bbb4b690bfbbc260bad3b5;
// music[695] = 256'hc6b174b36abda0c227c1aebe3dbb52be98bf7bbce0c332c677bd08ba44bf48c5;
// music[696] = 256'h98c332c788ca45c971cf3fc8b7bebfc692c94fcaf3cd4eceffd051d0b6ce86d2;
// music[697] = 256'h02d491d881dfaadcb1dbc4dc53d50cd57cdbb4d932d519d885e0f0e464e32ae0;
// music[698] = 256'h58e24ee5b9dd44da66e278e772e77ae797e9d5ea15e7c2e111dfbcdb69dc99e5;
// music[699] = 256'ha9e8bae57fe416e645eed1ea9fe5d2f3bffdcf03f80af405effe78fd44051b0b;
// music[700] = 256'ha006cd094d0cba07b408cd060405770811040c00bd023005210f890fd203ba10;
// music[701] = 256'h9e200020a122561ede1b11219d22fc27a82730296e2f88296a25b124fb23c625;
// music[702] = 256'hc6244f2a492ced22f5204224ae1ebf19fb1d071fc51f4c222e1f3b20b81f0b1a;
// music[703] = 256'h221b7e220e27d21e2a17bd17a41579140917121b891b211e8322421cf61cff1c;
// music[704] = 256'h0314f1194917460776086d088a01d0037b0186fb62fdf1fe24048608a9074508;
// music[705] = 256'h4f021f016b008aee38df2bd8dcded8ea8aeb32f1b7f116ee47f064e971e938ed;
// music[706] = 256'h97e983edabf159ee94e73ae118de4adc78dbb6dd44e1d7de14e2adeaeae0f6d8;
// music[707] = 256'h56e477e97ce804f3e5ff040282fde3fca501450255fc25f881f861f6f2f124f3;
// music[708] = 256'h1cef48e7a7e85debd4f265f8abf85801f3fd40f5d3fa570271075b036c024f09;
// music[709] = 256'hfa0693071d0ac60ad30df70f121604195019e9196e17491bda1dad1df520b520;
// music[710] = 256'h1820db20c921c62447295229702368267e2c392a2a2bb72cb72b552e722d2d2c;
// music[711] = 256'hf6325334562dc42daf31e732ce33c02c44289b2ece2d242ce32fb52b2d2a392d;
// music[712] = 256'h172aa827c328182de12d5329f3287625b8221127df28bb2c1d2e782647231225;
// music[713] = 256'hf823fc25bf2b13260b1d541eb61f582449264e1fd720c91e571cfa2d733a5c39;
// music[714] = 256'h003a233a3f395f38b738d334172dd52b71294928df2c432c352b012cca30a236;
// music[715] = 256'h2a31ab2f6e33642edb27d923822906310d2bcc2393208f2458322b347129c824;
// music[716] = 256'h45233924e523cb16d512d51bf81ae51b7d204a1fc31edb1f0b21f819b018bf1e;
// music[717] = 256'h260c04fa86fc73f9fcf669f8f2f581f6f8f5baf158ed19e82be4e2e048e09ae5;
// music[718] = 256'h84e27fd9e1db64db62d315d394d200ce62d03dd318cf0ed0b2ce17c612c9c5c8;
// music[719] = 256'h6fc0cec476c807c469be66bd20c261c083bfcac2bac1ecc2fec2a9c230c663c4;
// music[720] = 256'h33be3cba32bb92be1cbf7bbf63bf4fbdfdc02bc9b6cab8c935c979c248c02cc4;
// music[721] = 256'h2cc78dcee7cdddc975cd2cc882c7ebcfdbd010d31dd25dd074d0ebc8c0c9a5d0;
// music[722] = 256'h52d2e8d408d861d958d335d7efeac0f048ee07f097ec9deb13f2b3f88ffaa2f8;
// music[723] = 256'h9bf5c8f15defc3f03ff7d6fdcdfeebfe2dfe75fa69f77bf6c8fbd9ff66fbcffc;
// music[724] = 256'hfcfcccf5bbfa27030c05730365fae6f6ebf9c9fafbfc8ffadbf761fbb6fd5afe;
// music[725] = 256'hf9fee7ff2ffe73fb41fd94fc87f9daf8f5fb5d0344ffe0f45bf52ef6e7f42af4;
// music[726] = 256'h33f8cd00f0fdc4fbc1fc1cfbf701060072fc7601ea01c510a21cf916431ab319;
// music[727] = 256'h6e15a5198d19121a931cd21be61d0f1ffc1aa419bf1a2017c916311b041aef1c;
// music[728] = 256'h6b22051042f915fdcb005afcc500ce01b2004202c7fe12011308f1012afb22ff;
// music[729] = 256'h85febafe2100d8fb3402780404018c071c0433ff8cfc48f7920323048cf09be9;
// music[730] = 256'h43e50ae28de3acdfbfe433edd0e9d5e632e5c7e4dfe982e84ee5b8e9f1eb1be8;
// music[731] = 256'hbbe1c9dcd9ddd0e333ea4aed83eed3f2d6f3f6e92fe459e7d1eb0bf410f500f0;
// music[732] = 256'h35ed94e099d517d968dff0e13ee438eca6f168eaa4dd91db8be75af1bdf64af9;
// music[733] = 256'h0df82fff370611046103a2ff75fa9dfb68f5e8eb00ee99f151f322f7c7f867f4;
// music[734] = 256'h14eff2f279f34df3b8fbfcf792f50800a0051509ee07d10400046b03c106d80b;
// music[735] = 256'he11273127010d315321493182921b0245627191d2c194d1f191f70269b29fe24;
// music[736] = 256'h6329b02cac2a602d1230d52c242df02ca029602d24308b3418395a314a2ec932;
// music[737] = 256'h22310a2df02abe2a622b522db52fb42f3d2efe2b31299429142f9c311e313231;
// music[738] = 256'h142d7d29af24a2205d29e62dfc28c429552b632deb2af41fa721742ae8297129;
// music[739] = 256'h3c262c209e24032a35256323ac27c824a328ed38a23dcd395939d63d5f404938;
// music[740] = 256'hb037b0366c2dd1312734b22eab2dba2c05302231b5304c3396344c35582ec32c;
// music[741] = 256'hbc33622eeb28302abe28c3271f28db2cbb31932e182b5a297122821c091ec51f;
// music[742] = 256'h2a1b5017b91a691c741b721e361f7a1f2920691de21f6c20121189008bfca1fa;
// music[743] = 256'h37f60bf602f8bbf6d7ef24ed34f251f1d6ef2aee4ce512e580e50bdd46de6ce2;
// music[744] = 256'h36de36de73e081dbfdd799d716d2f4cd2cd032d3bfcf50c7c8c9e3cd46c594c3;
// music[745] = 256'hbcc616c34dc064bcf5c2add4e5dce5df11dec8d940d955d4e3d60cddead6d8d3;
// music[746] = 256'h99d640db6fdfa4d75bd36add6ade8bd69ad892dd5be246e619e0ebdde1df7cdb;
// music[747] = 256'h24ddefde6fdbd8db41e047e59ce29ce1ace6fee4efe5aae7cce7daec7bebf5eb;
// music[748] = 256'ha3eda5e5b5e23ce574e9c8e89de33aecb1f010ecc6ee8bed9aee78f2b0ea6be7;
// music[749] = 256'h0eefc8efa3eaebed09efbde7d5e960f33ef59af17af259f23bed3bedc5ee2df3;
// music[750] = 256'h2bf64ef086f1fff183eddfedd7ed7ff4e1f877f7b8f998f4d3f256f596f450f9;
// music[751] = 256'h2aed39d6b0d79cdc2bd6b6d6c1d974d78bd46cd9ede129ddd8da37de24db1fe0;
// music[752] = 256'hdcdf91da36dfbcde38e05be042e616fa1bfc1ffbb8ff7efa2ffbf8f8b2f408f9;
// music[753] = 256'hc4f9e6f7c3f92cfec1fc49f8aef833facafd03fd3af9f9fd0c03c2000ffea100;
// music[754] = 256'hc902b1038d02d6fb9cfa78fe550156045d0076fb77fd2f0092ff3efe45fe55fd;
// music[755] = 256'h58ffc100eefaa5f7f8fa1a05e2097ffea3f976f980ee29e6b1e2dbe6b8eb4de5;
// music[756] = 256'ha7e551e866e842ec41e6d4e2a5e2e3dff6e820eca3e89fe6a8ded8e1cae79ae5;
// music[757] = 256'h0becd8f196ec8dedc8f23bedb8e89be6ace690f099ed56e7c6e8acdf07db1bdc;
// music[758] = 256'h22dd72e0e8dd83e345e7c7da48d82be5a8ee4ff456f967f9dffe2b04ddfd40fe;
// music[759] = 256'h3cff34f94dfa35fca9f79ff2ddf444f63af555f565ef49f183f5f7f4b9fcc2fb;
// music[760] = 256'h62f8a2fa2bfaf0ffb202640348055505800b180c390fdf159e102513401ad416;
// music[761] = 256'ha513a0150f1a021bfc1c8f213423af25e323aa24692f5a302b29cd291b2e5c2e;
// music[762] = 256'h582a2a2c5332b53116337137dc340b35293894340d354f39e035662f082ba72f;
// music[763] = 256'h92375032d52cf02d4b2d732f9330e03149372b38423661333030843270356e31;
// music[764] = 256'hf0296327a12af42a05262523d024782ac02e402ad5289f2a7c2535246425fb25;
// music[765] = 256'hbf2569205b225f264c2b59378d37ad34ec38b2398a3a123751338f352a32bd2e;
// music[766] = 256'hc4305f317a30132f922fe431ad33be36e8358e30df2fe630b12ef42ccc2a2b28;
// music[767] = 256'h4f29bb29c32880320337842afe282f29ed201928092b0124a62630276c253722;
// music[768] = 256'h15204d246a1f74254a3b4c3f113fcd38f61f4b151017c318031ada1089102d16;
// music[769] = 256'hc211c911710d69065309b0058dfd3affcd0269fe40fbd1fd82f8c9f03df3b1f6;
// music[770] = 256'h62f1baebb1ea02e66de585ec50ec46e659e31be426e472dfb3d930da08deaedd;
// music[771] = 256'h67de03dbead21dd5fbd6a1d53edafedbc6d87bd4f1d3a0d426d60adbe6d690cf;
// music[772] = 256'hc0d2d1d6b0d239d093d4b7cfa5cc6cd461d681d80ed9afd6bbd8cad403d39ad8;
// music[773] = 256'hb7dc98dc5cd704d639d94ed96fd825dca7e026dfb5e0f4e24fde98e039e5c8d8;
// music[774] = 256'h4cc82bc662c653c8b7ce7dca00ca69d0e5cc40cd4dced8cacccfc3d0abcde0d2;
// music[775] = 256'ha2d41cd372d392d09dd3c2d9dbd868d858d677d4f9d57ed4b2d35bd336d5bfd6;
// music[776] = 256'h1dd243d4c8d9eddcb5e087dfb8dff1e241e32fe009deb2e1b1ddcdd503dbd0e0;
// music[777] = 256'h49df0ce084e1e0dee8df09e241e068e240e094dee7e493e30ee4d9e344dc2cde;
// music[778] = 256'h91dd7ae01cf2dff804fb43020802b3fe9bfcaafb19fea2ff41fb98f8bffd7201;
// music[779] = 256'h85039802a1f933f77efe0f023100470090feb7f888fde90299fd2bfe3f006d02;
// music[780] = 256'hfd03effbe7fc9f037c02a902a8ff88faaafb5302a906730386046005c800c000;
// music[781] = 256'h2f006d0211063403b302cdf969ea62e777e55fe6e7ebcfe7c3e9b2ef0ee893e6;
// music[782] = 256'h7feb27e7b4e798eb0fe813eb6ff0aae7d9e20dec85ee11ed81f1a6f27df3faf4;
// music[783] = 256'h3bf2a0ee6fe9b4ead8f3f3f54df0cfe91de6a9e299dd68de52e514ebaae881e6;
// music[784] = 256'hc8e7a3e057e0f2e93bf012f9e3fe19025203fc025908a4040501fa033501e100;
// music[785] = 256'h14fa22f4b5f679f140f462f735f1e2f64afd56fc8cfbb1fa74fb75fb2afdd9ff;
// music[786] = 256'h2101fe02a904c309fe0a910507094e100f119e11301426159114161adc200620;
// music[787] = 256'h51231426a0224227a02cba2d1c2e7d2af62b102d07298d2bc82dc52def325837;
// music[788] = 256'h00389e35c7317d325c3564331e320a352f36b538ff3b8f3809358a335f2fbd2f;
// music[789] = 256'h1235b2385a3953370538933802341331fa34363bdd369e333b391532e72d1d33;
// music[790] = 256'he7301f338f326a30eb31be2bd12ba32c8429f22c832b7328b8278126d623db27;
// music[791] = 256'h12390d3e0f416052df56ef555556c3528f54cc51864c864be248d44b14518a4e;
// music[792] = 256'h8e4a554c334f324f8a5067503b4b9547d8474748a647c24548414c3fa046894f;
// music[793] = 256'hf24eac4665403040b63e053c6f3d3d3c09374537fb3b483b5139813b123abc39;
// music[794] = 256'hef382034da33a7278d167a1644136a0e4f0f5a0bdc0aa40adf05eb02feff80fd;
// music[795] = 256'h49fc3ffc1efd0cfdd0f70aee3fe94ee855e808e8a2e454e4a4e6b2e53ee078dc;
// music[796] = 256'h08dfc2df0fdf44db04d6b7d7b0d44cd37dd71dd241d1bdd43dd49cd3abc47cb3;
// music[797] = 256'h6eb14fb3e0b546b532b1e7b108b49cb3c7b114b0fdaf3fb185b20cb4e1b143ad;
// music[798] = 256'he1b1efb6c9b253b3edb64fb62eb6e8b53db8d9bdb6bd94bba3bb77b922be09c2;
// music[799] = 256'hf7ba6abeb0c4b5c1acc287c1d2c11cc42fc418ca0fc988c5b6c8bec7b7c8d0ca;
// music[800] = 256'h14cc48ccbac7f7c9accefcccfbcc2dd0bed212d299d18ed2dcd1f5d1dad389d4;
// music[801] = 256'h6fd5a5d90bdaccd89fdc86d930d5efd87dda3adb53dc06dd41dedadbb1d8f6d7;
// music[802] = 256'hefdb56de4ed99adaeadf16ddeadadedd68ded6db67db09dfa3e0cddcd7dc65e0;
// music[803] = 256'hecdfece0d6df2fdf6ce5ffe30fdf83df20df6edf7be1fee4c0e29ae651fa99fe;
// music[804] = 256'he1f9dffc56f917f9ccfbb3fccd00c4fee0fc3afe28fe8bff29ff6ffdc2fc50ff;
// music[805] = 256'hd30186fef9fc3efd3ffd11009efe4cfb2200770484020b036c045204d1042e02;
// music[806] = 256'h50029205110451036f03a6ffb4fe1704fc070e0624041003c8008cff87fee301;
// music[807] = 256'h430417f514e81aece4ea08e8ece98be981ec22ec7aea3aeb89e827ea2aec05ee;
// music[808] = 256'hb8f051ed5bea53e5fee2afe8aeeb0fee77eea1ef0ff392f1b2f23af12eea8dec;
// music[809] = 256'hddf082eddcebabebabe6f0e33ee218dfcbe075e1e7e59cf046ea62dd9fe2c7ea;
// music[810] = 256'he5ef53f848faebfd7204ff039205150346fd66ff27fdf5f6c9f5a2f740f577f0;
// music[811] = 256'h2df2b1f3edf33cf4d4f25af5d9f7dffa0bfd0200bc04fe00e9019d078608af0c;
// music[812] = 256'hd40d5c0f38125c11ee13cb16211a941a301b9e22f82524283a290728912a8d29;
// music[813] = 256'h2c2b6e3015314632d7345b367e35ef34bf347935613a9c38543541375f38863c;
// music[814] = 256'hda3a713eb9514658a055e3563958185bbd572455a955c5521c54455354501e50;
// music[815] = 256'hb64e18522c53ed4ecc4e794e7a4d1a4e914ef54fc94f944ec64ea14c47492448;
// music[816] = 256'hdf477a474b449844b5482444fa41e9434040e63fc63e02463357365779524d54;
// music[817] = 256'h1954a854e552d9533c53f14c4c4de74a5d46fa47f74553439c45fe49034c2e4a;
// music[818] = 256'hd846e4410842ef428f3f4f42ee410b3c2c3afb37dc3d58462542b23c9839e735;
// music[819] = 256'h89345a33f833ab353f347b313432e33217314c30402d302daf2f7626f213a3fe;
// music[820] = 256'h6bf20ef3f3efaaeca8ef25f029eca6e871e8fce59ae1aedd6adb35dc04d98fd8;
// music[821] = 256'hfad808d17cd093d286cc9cc90fca0fcac1c64cc450c60bc436c220c291bf02c1;
// music[822] = 256'h1dbf24baa9bcafbea4bc42bab0b764b6beb5d2b6a4b763b794b882b6b0b2b5b1;
// music[823] = 256'h78b33fb71fb856b7a9b4b5b03cb4ecb636b523b8a3b628b38eb8d9bafeb798b8;
// music[824] = 256'hf4b86ab8f2b61ab7c4baa6b987bb2cc22abfcebc71bfcbbe76c087c2b9c234c3;
// music[825] = 256'h72c2a0c311c5bbc41ac41bc42ec7bcc67bc348c7d3c98bc9d8cd3dce1acc6dcf;
// music[826] = 256'hc6d11cd101d3fcd510d6a7d7afd800d601d8f9d811d5e4d495d58ad85add0fde;
// music[827] = 256'he6dc26db49dbd6dbb9db51df39e132df80df06e2a5e079dc8adb19db1ad9c4d9;
// music[828] = 256'h03dfebe013dd1ce0a5e4afe2e5e394e633e736e6d1e424e787e6afe2e5e374e4;
// music[829] = 256'hc6e1ffe3f7e746e6f1e27ae2ece3dcdf7fdc54eb6dfac5f9d5fb59ff9cfd10fe;
// music[830] = 256'h2efd2cfe6503000134fda8fdf9fc5a012c0334fe64ffd7003201730245017c04;
// music[831] = 256'h0e060d03ef016402af040602defffd0328032f039a07ed05b001d70157039d04;
// music[832] = 256'h1b07ca068b042505ea066d070a0633077e082b04ba025f07fe021df1dee8b5ed;
// music[833] = 256'h3eec2fec46efdeed97eea9ed81ea0beb58ee00ef18ebf7ecfef0baef91eb98e5;
// music[834] = 256'h98e858ef52eec7efdaf2a2f285f1ecef64f1ceee5de9cff1c8f931f210ed4deb;
// music[835] = 256'hf7e768eafde733e3ebe7abeb09ef08f2ebe952e51fedc7f3d9f9f400f805720b;
// music[836] = 256'h090cb2086109610bd308d602110178ff6cfb11fa33f952fc65fc58f9e2fcbefa;
// music[837] = 256'h78039c18601d66201822ca1fd226ea26b226242ca62b102ed130ed321e378835;
// music[838] = 256'h9934f237dd39ec39203c07409b3e503e2645f448a3488348684794492f4e884e;
// music[839] = 256'had4e0952085488534d513b5022547f56d852eb507a51ea5280558553ba53dc57;
// music[840] = 256'h62569d561d57f05465580b583b532b542a55d551ec4ca94bc34bd248824ab94e;
// music[841] = 256'h7d4c5a4a834ba3496c4733485d48ad47fe479349894788412d3d223b613ea83f;
// music[842] = 256'hd63a493bf9397c36f33720356a370c479050124ca34be74c393eca30932de628;
// music[843] = 256'h0729d82bdf29b4255b247525a825cc25c225042afb2bd82768296d2788254428;
// music[844] = 256'hef230721781ea41ce51e6a20642877289621fb245b22671b4a1dc11dbf196d17;
// music[845] = 256'hd218381bc11a021bde1c76188216dc19cf17b816760c52f9d0f4f5f270ef9af1;
// music[846] = 256'hbfee2fed0ceea2e74ee366e4bde005df38e255dde5d6f5d5f1d353d3b6d3fbd0;
// music[847] = 256'hc8cc63cbecca98c84cc8c6c8c0c6e2c2c8c0c5c183c02ebed5bb82b902ba09bd;
// music[848] = 256'hffbde1ba68bbd7baccb58fb641b8c6ba18bbdcb76cbaafb8ffb5d3b785b7e5b9;
// music[849] = 256'h92b750b69dbacdb66ab4c1b668b749b6e5b39ab76cb9fdb529b9babbb3b9a0b9;
// music[850] = 256'h08b849b81bbdecbdf4bc86bd52bf67c4ccc405c2b6c502c832c400c2a0c101c1;
// music[851] = 256'h28c3c5c31ec544ca09caf8ca40cd52ca4bce9bd341d4d2d5a6d520d694d65ad5;
// music[852] = 256'h3ad63ad846d797d409d781d920dac1d99ed6c9d9f7db03d9f5dbc4dc30db9cdf;
// music[853] = 256'hb5e29ddf9cdfe0e1ecde00e168e464e1f4e138e33ae3c8e063dc2adf25e21ae2;
// music[854] = 256'h95e2c6e244e37ce1e5e289e72ee748e640e6aae46ee437e3bae0ade355e6f8e3;
// music[855] = 256'h63e1f9defae10ce621e95df82a0397ff8dff47ffeffb6dffbc01fcfe36013a03;
// music[856] = 256'h2e02f203610083fdcf01d302ff015b0066ffd5027004910345022c024403c502;
// music[857] = 256'hef006f00e902e503b504b4076a050a036e058703d001d006a6061e020605490a;
// music[858] = 256'hd50bcd0a0b0892078e0a280afc08bf0c340234f118f240f011ec93f0d9f09cf2;
// music[859] = 256'hfef241f173f481f470f309f400f613f76af5b2f3d9efc6ef25f303f3b0f44301;
// music[860] = 256'he614bd1aea18401b421770123f1380176b17dd1042117e0d6d042c078c082504;
// music[861] = 256'h8306c00a2c0ef70db30320028a0f0b1540199b2249243925de28042866235d1f;
// music[862] = 256'h0b1e021dc91a8a164414521533156514ab130616af188b1583148e182b1c901c;
// music[863] = 256'ha61a311b7e1dcd20ea2543282d29982c8e301f3219311d338235aa315232e136;
// music[864] = 256'h2635433315358a3a513cfe39354120467e43db45554750475047fe443c452f46;
// music[865] = 256'h7746dc472248f646f7457746f9494d4b0e466a46bb472c39772a1528ac29b82c;
// music[866] = 256'h1e2dbe2b782d0f2f5b309b2f8a2aef2a222eac2a38286026a1230e27072a8e29;
// music[867] = 256'h0e28b2251a26f4251a237c24f228e9264a249d263d224a1c0d1ae218011c371c;
// music[868] = 256'h751db91e701f9d2ff837a530fb31553344321c31ca2c0e2c212b7d29ac282f26;
// music[869] = 256'hb925fe28b12a3b268827482da02946252c247822ef2205242623b921ab22481f;
// music[870] = 256'hd81ca9267b2d6029d422131e641c5c1a3f1813189518c3170019491cc1197719;
// music[871] = 256'h521ada1533177c167613f412870541fadbf925f46ff1f6f280ef63eccbecfcec;
// music[872] = 256'hace875e528e597e1abdeebda87d7f6d827d7d9d6a0d70cd29acf5ace4ecac8c9;
// music[873] = 256'h82cc85cbd5c4a0c48dc74ac5d3c2b0bff6c027c2acbe92bfc7bdd6ba93bb11ba;
// music[874] = 256'hf6b720b7b8b958ba9fb707b9b5b849b875b914b64db616bbf2b6b0b030b415b6;
// music[875] = 256'h00b5f1b638b6b1b78dba87b932b949bbe3bd9bbb17ba91bc80bb50bc64be16bd;
// music[876] = 256'h18bc23bdc1c0ccc16fc153c2a1c1d7c253c3abc23ec722ca10c873c73ac648c5;
// music[877] = 256'h58c821c857c955cf45cf10d1dbd3dace2cd06dd46cd2add1e1d2e2d4acd4c7d2;
// music[878] = 256'h60d4fbd64bd859d7a7d7b2d942d81dd86edad1db64dbf6d94adcc9dd0edc2edc;
// music[879] = 256'ha7dd9ee18ce321e085dfe9e379e548e291e2b9e5b5e610e633e3a4e3f6e66be6;
// music[880] = 256'h58e5fae5abe66de8fdeae0e828e35be1e5e3dfe5eee26ae118e20ae20de715e7;
// music[881] = 256'h2bed8800d0035b015b05c1048d060906a0038203c10181038a052c03f2000104;
// music[882] = 256'h060a7d0ccb0b59089607be09e409c509e10be30d660ac70cdc0f890a9c186a2a;
// music[883] = 256'he628e7272529cd2c6e2cfb28ba2d4b2b9a28f72b742bf42d472d092ad8292429;
// music[884] = 256'h8129fe276d2ab2286316e60e8a142310660c0e0d140b370c480b300bac0f0f0f;
// music[885] = 256'h250ffb0f8a0e1213c4157811390c530b670e9d0e60101b147213a31443189517;
// music[886] = 256'hf81322125712fb138c12ae0cda094607010527066605a906e2070a0b3511e606;
// music[887] = 256'h51fa5000dc071f0e4219771f3d201720811e281f8f1d8c163a151a14da0f8d10;
// music[888] = 256'he20e600b0e0af907e3066807f90a6c0a10094f0cd40065f06fef72f28cf7b3fb;
// music[889] = 256'h98f8a3f8d3fb7bfff7044c068407310ac10bb00fe30f7b1188168a12b5121019;
// music[890] = 256'hc4194b1b071df31fb921b4205f24c3257226f027c225f32687278b27fd28a128;
// music[891] = 256'hf02a342c8d2c452f052f162d5f2c0a2c632ba32c362c672a4b2fbc31ad2db12d;
// music[892] = 256'h472f872e072e2d2db22bf82e283021292a29542d952a6a284327d325ab255c27;
// music[893] = 256'h42296b26d123e224d5251824a8201b204c20f91d301d411f251cbf196828a334;
// music[894] = 256'hd1312c32f631a13233371731be2e4434d62e9a2a162e7e2ce2299b2aa72aae2a;
// music[895] = 256'h152e6131082fd32cec2b41290e2950275724a0249e2221200c24f82a802a8225;
// music[896] = 256'h9924c1215b20e921181f0e1f801dc218a11c511f0d1e8b1e301bf61ac41b8317;
// music[897] = 256'hea187d12cfff44f9ebfac8f915f535ed29ed15f0d1ecafe748e336e268e3b9e3;
// music[898] = 256'h47e122dd91da31da8eda39d61ad445d529d0fecf20d1cdcbe1c8b8c69ac9c9c9;
// music[899] = 256'h1dc3eac5fbc4c4bf0fc396c169c042c38dbf73bdefbda5bc91bc1cbbb1ba75ba;
// music[900] = 256'h5fb795b9f7ba0eb644b5ceb5bdb461b50eb502b5f2b532b7b0b79bb71cba76bb;
// music[901] = 256'h99bbaabc1cbc26bdddbc34b9d3b867b956bb96bf5cc0fdc065c293c2e6c21ec1;
// music[902] = 256'heac131c512c4cec457c865c8f5c78bc935cbffcac2ca60ce77d0c6cc3acc1ad1;
// music[903] = 256'hd0d3bbd4b9d50cd5c3d30ad480d511d6acd5bed68fd9fcda4edba4db20d952d7;
// music[904] = 256'he8d8f3da39da2ed8bcdb42df01e18de43ee225e3cfe6b0e224e3f4e870eb8dea;
// music[905] = 256'hcbebc5eed3ea41e9a2ec74edd1ec5eeb15edfaea2ceb72f1b0ec52f3dd07680a;
// music[906] = 256'hc60685076208670994075f08480ab6077e054e061e07a80b52191a22da1fb91f;
// music[907] = 256'h1f226222e02369266125eb231025d4239d24b327422545216b206b24f2269722;
// music[908] = 256'hd6222424cf21ec2540276424672620265f26b0279125e825672563267729a826;
// music[909] = 256'h17268c26042511273325dd23cd2656245023bb26b625b224862548236b253322;
// music[910] = 256'h750e6108cf0fd6097a040507d9075a07c406a206e9037503ae043203d9067e0a;
// music[911] = 256'h6807d100e6fb87fd03008d025005a007d708acfbc4eb8be99ae545e327ed1af1;
// music[912] = 256'h06eb93e82ee583de19dc42d977d8bcdce6df54e77fea9fdef5da1ce481e629ec;
// music[913] = 256'ha0f8cbf932f991ff6601b100a2ffe9fa88f7fbf54ff25cefa4ef72ee2bedffee;
// music[914] = 256'h3af0d4efd7ec5eed7af204f107f2dcf88ef849f9ddfeafff3bffb300f7ffc502;
// music[915] = 256'h5f08d205b505a70b730d5512ab13570fc912f0161a19511a8c1a071d411d0b21;
// music[916] = 256'h8b24a02341277b25452362282827b5258a2ae52c7f2bef2adf2b272ddf2f302e;
// music[917] = 256'he42b3b2fd12f8c2e2c2d072dc930ce2fa32e8f318a317131d331212ff32e0933;
// music[918] = 256'hf430002e3632ee2fd92b352d452b6a2bd42b8a29822aee2ac429ae277727242a;
// music[919] = 256'h8927a4232e235921821fc81ee01dd41d1c1ced1f6931f33ab1333030c7325237;
// music[920] = 256'h3e37ae2f282de42a582aea2d262b5e2bb22be729272db32d0c328c31a129232d;
// music[921] = 256'h642c15279b28bf26a527b42a062998268128bb2ecf2d23292527b122eb20d220;
// music[922] = 256'hc21ffd1f3b1cd2182c1a71194e19081c3a1aeb176d1a911c361aeb0e1e00acfb;
// music[923] = 256'hcefc74f770f286f3b8f189ef23ee2de824e785e830e547e2a5dea4dcecda2ad7;
// music[924] = 256'h8cd691d5cad232d244d3b1d15eccbcc8e9c60cc783c7b9c47fc2c0c162c3d2c4;
// music[925] = 256'hf6c079bf7fc1dfbf44bc6dbb90be0fbf3fbbeebba9bb7ab716ba33bc45b9bdb8;
// music[926] = 256'hbeb829bb8dbaccb533b84ab92bb789b93eb9e5b569b5eeb8acbb88ba10ba02b9;
// music[927] = 256'h99b7f2b9bfbb1bbdecbfa6bf93beb8bd2bbc6bc00fc7cdc99bc81dc547c77fcb;
// music[928] = 256'h4ec9dbc9dccf31d17fd160d414d20cd137d30fd4efd5bdd5dee290f57df4f2f5;
// music[929] = 256'h94f93df4aef660f77ef49af7a1f936f862f8a1fb21fc99fc79fd1efbd2fe3802;
// music[930] = 256'h01fe45fecc0242019dfe8fff1b006802c2049205d4065005a10578064506b607;
// music[931] = 256'h7007f606a505e604f904540354044403bb02f905690888095d068a0414045403;
// music[932] = 256'h78068c06b606c10558049407aa03040722192920321e7b1f2a20651ec21c841d;
// music[933] = 256'h4e1ec51da01dab1c2d1cd51c4c1aae17cc174d183e19a91726178d192c1a0e1a;
// music[934] = 256'hf918261a441a2c18c2195119a01c2b1cc20922fdeafcd0fc65fde3fde6fe0cff;
// music[935] = 256'h41fec6fdd7fc82fdd4fd2bfd37fc35fc3ffdf0fe85fdb3ef46e287e31de571e2;
// music[936] = 256'h0de3e1e451e590e5bde5c9e5ade53fe484e351e5c0e7c5e9d0e7c5e037de73e3;
// music[937] = 256'h8ce520e8ddef83f001ef87ef68ec90ece8ea58e9e0eff6edaae6dae607e2fdda;
// music[938] = 256'hf8db33dbbed931dda7e082e6dfe4a8d72ad997e571e9a7ef41f764f9aefc26fe;
// music[939] = 256'h9bfd91fcbaf8d1f6a9f5c2f2ddefd4ed41eea9ed08ec0eec05ed0aef33eec4ed;
// music[940] = 256'h18f14ff34ff4b2f3d3f575fad2fac1fca0ff41009902e9045d08ec0b1f0d1d0f;
// music[941] = 256'h7e1056100112dd14e1151d18d31c621eef1ef7204c223024ee24e32467279c28;
// music[942] = 256'h97272628ac296b2bb42bd629cf2ab52c342d082fc42eec2c002c9d2bb52c472d;
// music[943] = 256'h4e2f2f30f92dd42e0b2e232da52f4d2fc42e532e8d2e6330be2f7930d02f892c;
// music[944] = 256'h1d2d072ee02c612c4c2db72d572c152b6f29de2733270226af23bb235a241b21;
// music[945] = 256'h3621452207201c204b1e15244933c2372e3548353137c837e2347d3458330330;
// music[946] = 256'h1e310931442dc02b8b2c1e2c2f2be52dfd30b52ea62cd92c882aa6299f292828;
// music[947] = 256'hec27a22575233f248c29c32fc02b4427f0268521071fde1fc01e661e4a1eb61d;
// music[948] = 256'h461c7f1b901b211b421c4a1c631af21b9c190e0920fbfdf9cdf753f5f3f466f1;
// music[949] = 256'h40ef04ef64ed02ebbbe750e39be122e116dd7fdabcd99ad73ad745d625d3ead0;
// music[950] = 256'heacff4cc97cad9cb43ca48c6ddc517c993caf8c530c4bfc66ac677c5b1c4b7c3;
// music[951] = 256'h9bc33dc3c1c2a5c2aec136c0e7bfdabe94bf06bffbbc5fcb57ddafdd78dbfedb;
// music[952] = 256'h5adc0fde63dcd1dbe1dc77dc3cdd13dd9eddf8dec0dda8de1be0bdded0de3cdf;
// music[953] = 256'h7fdf69e0e2e08ce2e3e19ee11ae5efe3e4e2d6e651e7e2e621e8f5e6c5e612e9;
// music[954] = 256'h63e90cea0dedc2ed36eeafef4defdbf12ff598f337f2a9f22ef3d4f48ef5dbf4;
// music[955] = 256'hc1f498f515f7e7f709f81df9fef930f9bef7d1f773f9c3f979f93bfb79fc0afd;
// music[956] = 256'h81ffecfedefb82fdc6fdf8fb71fe62fd05fa1cfb89fc9efcd4f931f969fc97fb;
// music[957] = 256'ha7fbdafca1fce3fd31fba7fbddfb00ea35db24dd0ddc54dae3db93db2adfdadf;
// music[958] = 256'hb9ddd5de6fdd4be758f980fc65fbecfc6afb4dfb9cfb0efc4dfd3afda6fcddfc;
// music[959] = 256'h41fea4fefdfdc5fcb5fb90fc84fe0700e8fe71fdecfeb70012004fff6e031d05;
// music[960] = 256'h4602f903ea039701800179012e03660116009102440114034c058a02e9003000;
// music[961] = 256'h230219022c00900197ffd0007afe0dede9e4b9e7bde57ee533e5f3e321e5f3e4;
// music[962] = 256'h5ae565e552e5bbe7c6e74ce671e8f4eb9ce874e13ce305e870e8d8ead5eca1ed;
// music[963] = 256'hcdef22ef05ee80ece1e821ecc6f14ced19e6c0e367e1b6de03ded8deeae0bce3;
// music[964] = 256'h5be9a0ec12e3aedbf1e3e1eae2eee9f79afde6004104cb037a01ebffbffe02fc;
// music[965] = 256'h88f89af51af4a0f4eaf3d8f2fcf147f19af14fef10eecaf19bf45bf5c6f709fb;
// music[966] = 256'hf6fb48fc6efd53ffab0262067c0901092e08ca0bb90df50da21088149e179e18;
// music[967] = 256'hfd198d1bbd1cfd1eb421e3246127b029cf2a5729462a582d9b2d9a2b582c952e;
// music[968] = 256'h042eb22edf2f072fd82f0a30702f9630fd30f32f3c2fea2f5d3192319831a432;
// music[969] = 256'h07323a31ce32d132e9326034ad32fb304e309d2d9b2d603048304c2e632e6030;
// music[970] = 256'h732f342c242c5c2b032a6d2ba22a212a68282923bd2274221d20be202b21a01f;
// music[971] = 256'h36204a2cad384d3786355c367b38493a6a35d33425352331f230c52f1f2f292f;
// music[972] = 256'hb82cf02cac2dfc2f7d31cf2e592dc52b182a5729fc282c292727b22568247425;
// music[973] = 256'h0f2d2e30032dae2b58295125dc238d237f2249220e2200224223b3236d23b522;
// music[974] = 256'heb22a62313244c25401dac0ac900070238fea6fbc40b5b1ab71706165d155211;
// music[975] = 256'h650e770a23093108e1055b045b003afeccfe6bfc4cf8bdf68ef555f1d1ef88f0;
// music[976] = 256'hd7ee8bec18eb5aeb53e981e6dfe5b6e488e4fae2e6e0f4df12ded1df82e08dde;
// music[977] = 256'h93dd01db70db57dc98d952daa5dcf2db15db89da1ed9a5da03dcf2d939dbf4dc;
// music[978] = 256'h59dc30dd11dc16db09dde7ddf0dc9bdc63dd51dd37ddf8ddc7ddaedc7cdc00dd;
// music[979] = 256'h54dc93dcb5de15e08fe0fee08ce0bddebade25e0bfe086e2fee364e4afe4d5e3;
// music[980] = 256'h1be37fe43be501e43eea71ebd6d74dcb35ce3dcdbcccbccd37cd42cecdcea5ce;
// music[981] = 256'hcfcee2cf4bd12ed145d021d002d1ced1dad225d4ebd571d7d3d896da47dac2da;
// music[982] = 256'h9bdc9cdc2add8cdd99dda4dc64dbcfdd2fdf4fde9fe03ce372e2e1e13fe257e1;
// music[983] = 256'h19e272e222e267e342e323e4b8e41be324e14adeffddcddebddf13dfb5e136f2;
// music[984] = 256'h47fd1dfb18fb6efa45f932f9b9f8d1f9e1f924fa25fa2dfa2afbb0fa2cfa1bfa;
// music[985] = 256'h52facafa4efb86fb80fa06fb19fcbcfc56fd05fdd6fc40fca8fcfdfd9efd87fd;
// music[986] = 256'h5afebbfe12fe5cfe80ff9cffd3ffe1ff0400710019007f001a0192000d00cfff;
// music[987] = 256'hcbffc60039f987ea21e802ebcbe815e9b2e865e8d1e800e8fbe8dae803e9c4e9;
// music[988] = 256'h78e9a7ead4ec57ede8e6d5e101e548e6f1e7aeecd5ed62ee35f076ef33ed3bea;
// music[989] = 256'h2be966ef50f279ec7ee998e629e2cbe01adf2bdf24e1cae237e793e7d8dd4adb;
// music[990] = 256'h69e604ed7df264fbe9fe2f02d3039602d5024c00e2fd5bfc3efaeef8c2f612f5;
// music[991] = 256'h1af469f3eef220f24bf2ddf220f453f560f6acf7adf8a8fa14fc75fdd6fffa01;
// music[992] = 256'h42054207bd07e909f80c960f4c11b6129914fe169e187c19351bf01bc11c7d1e;
// music[993] = 256'h2d1ff6217c250926de2655293d2bc02b9e2bee2b972c142d702dea2d9e2ed22e;
// music[994] = 256'h372e702e522fb92f6930ce30c33036315f310932b33283318d317232bf311832;
// music[995] = 256'h1932d5316532b4304a30a6310a31112f722d542e5c2e042e4530613170317530;
// music[996] = 256'h10306230e12e282feb2dd42a9c290329c428c12688260e271b2a8737363fc33c;
// music[997] = 256'h2a3c1b3de93e1c3e553bce3939398a373336164587563c55c05249531953b656;
// music[998] = 256'h345613531b52d550ab4ff54e854e524de54b2d4ad148784d5a534c505e4bfa49;
// music[999] = 256'h9b454d42c6413c3f053f5e3f573e3e3f173fd53ee13e9a3d693dde3bff3a9e3a;
// music[1000] = 256'hbf2e701f611cdb1b32186c16741449127e10bc0ea20cdc095608e00543035e01;
// music[1001] = 256'h97fe03fd0efbf3f83df798f42df27dedf5e957e9c5e7f4e6bbe50ae4f5e22ce1;
// music[1002] = 256'h44e074df52de00dd05dcc2daa7d73bd60dd68cd5e8d47fd3f8d213d206d22ed2;
// music[1003] = 256'ha6d178d2d3d0e6d238d024bb4dae03b1b3b001b1fdb10db25bb336b3c8b348b4;
// music[1004] = 256'h27b4f7b4fbb403b595b57cb656b7cab715b838b885b946bae6ba1abd56befebf;
// music[1005] = 256'h81c14ac1edc122c27bc2a5c300c4bac440c5e7c682c99ac92dc900c97bc9e5cb;
// music[1006] = 256'heecc7eccd7cc92cd03ce95ceffcfa4d0a5d069d1dad180d217d313d3d5d32dd4;
// music[1007] = 256'hfed3fbd456d727d94dd8c2d7cdd860d87dd8dcd918daefda2cdc54dcc7dcbcdc;
// music[1008] = 256'hccdbb6da55d97ad9cada5cdb33dc35dda3dd9cdd20de33df26dfe1df6ce1dce1;
// music[1009] = 256'hc5e20ce350e27ce117e15be2ede122e2b7e3f1e0c7e5fef401fbbff962fb9efb;
// music[1010] = 256'h38fbb2fb7efb82fc09fdf0fcb7fd81fdb3fdf7fd70fd37fe1dfeecfdf2fec8fe;
// music[1011] = 256'h5cff0f009cff550097003fffbffd0ffebfff18007f001a01b100e2000201e200;
// music[1012] = 256'h27015d01a5015e018d01cd01ff0079017001e000b2013500e7006e015af4ede6;
// music[1013] = 256'h80e71be90de826e97fe9d2e998ea99eafdea83eb85eb92eb59ecd6ed29f0cdee;
// music[1014] = 256'h6ce7a8e5abea45ecacee4ff268f23ff372f3d5f1efef04ecd9ecbaf26ef194eb;
// music[1015] = 256'h56e91ce610e23be138e04ee0e7e2f7e6c2ece7e7e7db74e08feb57efccf696fd;
// music[1016] = 256'heaffa803e1034202bf016cff92fd67fbcef8c9f770f670f57cf415f311f301f3;
// music[1017] = 256'h08f3ecf3c6f472f639f87bf9defa25fc17fe2e00c6025907b50ab60b430dbf0e;
// music[1018] = 256'hf40ff111651324158d17d918711b7a1f39212922aa232125fd27652a012b262c;
// music[1019] = 256'h122d362d582e352f9b2fc1314d338d330e363338ce37d937e2370e389838b438;
// music[1020] = 256'h7b39fe38af3877399138e7390539e838ec4a725c025b375a4a5b69575e56a354;
// music[1021] = 256'hd3522b54bb539853f3539b53f153ec528d5265521651465193502c501c50b64c;
// music[1022] = 256'h2e4be64a4a4975492d48b647a247bc44254cc8584a59fd561a58f858c45a3459;
// music[1023] = 256'h7a565656745401538c520651d6507450ef4eae4e2d51ae5317526350e64ff54d;
// music[1024] = 256'hd54c184a7d465d464445a542a3439749384d58489144fa42c63d073ce33a5e38;
// music[1025] = 256'h5e39ad388b3819387e3498356f3570332234fc30ab31142f6a1e4115b1141712;
// music[1026] = 256'hb710200def0c510716f011e27ae201df06dd10dce5d8cdd74cd5b8d284d145cf;
// music[1027] = 256'he6cd3eccf5c974c8dec601c6e9c4dac247c1d2bfb5be10be31bd4ebc45bb2bba;
// music[1028] = 256'h4bb9ccb8a2b878b85eb8ceb7f4b6f1b566b4f8b459b753b708b6c1b55cb5feb4;
// music[1029] = 256'h0bb5e5b4d4b4feb4f4b4b9b4b9b404b578b504b677b6c2b604b733b74fb7a8b7;
// music[1030] = 256'h1db897b828b947b995ba23be45c038c034c027c096c164c3b6c25fc2bac249c2;
// music[1031] = 256'ha1c2dcc22ec33fc48bc44bc5e2c5b7c57fc7a9c96dca2acbeecb86ccaeccf2cc;
// music[1032] = 256'h99cdfdcdf3ce96cf36d0c8d23fd400d4e5d4aed5f0d59ad62fd7c0d75fd8ded8;
// music[1033] = 256'h14d98cd95adac0daa0db92dc2ddd3edebbddb0dc5eddc7dd60dedadebddda8dd;
// music[1034] = 256'h9ade5cdf52e00de164e296e265e0eedfabe129e353e442e403e3e4e2a5e374e3;
// music[1035] = 256'he6e30ee5fae41de61fe622e526ef0ffd1bfe37fb67fcccfcaefd46feb5fdc9fe;
// music[1036] = 256'h7bfe30fcb7fbf1fc13fe9ffe61ff3e00b90074010d02950232037703eb03df03;
// music[1037] = 256'h9503f9032b04ad041305be04bf042a0448030303e302420344034f039c030103;
// music[1038] = 256'h4b03a1036203e203e702a302b5024c015e0337ff4df0d2e907ec5feb1ceb5aeb;
// music[1039] = 256'hfceaabeb6feb28eb95ebb3ebc4ebadeb1decf6ed7def5aebdae488e6ddeaa4eb;
// music[1040] = 256'h16effaf125f2a2f3e6f288f0a1ed53ea41ee50f302ef76eac3e823e4a3e150e1;
// music[1041] = 256'h7ae01ee4eee86aed41f007e6c6ddefe72ff01ff46dfd890126041d08a7060806;
// music[1042] = 256'h20052602d900acfdd7fc8afef0fc22fc6afb1dfa58fa07fa2ffb89fc78fdd6ff;
// music[1043] = 256'he60049043507c906a00ad30ac70c6a21d132463477365b383438753a953bcc3c;
// music[1044] = 256'ha23ee33faf41af42d7444d48c249a34ad84bc04cda4dcc4e5e4fd14f84505051;
// music[1045] = 256'h805196513952e2522f5438562356d054f6542055585595553f558f551055ba54;
// music[1046] = 256'h90555955b55567552b53bf52e15290520253005318539d51c94d774bd84ad14a;
// music[1047] = 256'h3b4b134b074bd04a104a264aaa4a40498a462346d645e643b243cf429f418e40;
// music[1048] = 256'hce3c4f3cf53adc39d8466a51424f1c4e4e4c9e4ca04e6e4b064b104a0248d548;
// music[1049] = 256'hf4458d476643bb2cca202d25c1271c29e9274d268925812264223b22db20be21;
// music[1050] = 256'h9e1ff91c9f205427b82740221d200e1dfa1704175615a314a115e2135314c414;
// music[1051] = 256'hef1304157414bd141b1480116812460a67f9a0f383f4d8f37af347f097ec28ea;
// music[1052] = 256'h22e7d7e4ade2f2e0bcde78db6cd9b7d7c5d592d387d1f5cfb5cd98cc7acb5ec9;
// music[1053] = 256'h5bc85ec6b9c40bc4a8c153c1bdc253c133bffebd88bc9bbb10bbdbb92fb9fcb8;
// music[1054] = 256'h26b842b744b660b5d7b404b473b3fdb28bb22eb3c2b355b32bb335b354b3ecb3;
// music[1055] = 256'h3fb4a3b4a0b56eb6c6b6c1b621b7d4b719b8bbb884b957ba76bc59bec6be10bf;
// music[1056] = 256'h55bf41bfaabfc5c0fac0dcc005c246c2c1c249c525c61ec6acc673c6ddc639c7;
// music[1057] = 256'h55c8ccca75cb88cb20cccacc0ccea3cd79cc27cddfcd49cedecf29d14cd11fd1;
// music[1058] = 256'h90d14ad388d4dad5d8d70fd78bd63cd8b9d896d952da90da5edbd9daa2db19dc;
// music[1059] = 256'h49daa7dab6d9aad8e3db0add62debedf00de0ce9e7fba9ffcdfc7ffdcafc7dfd;
// music[1060] = 256'hcefecbfe2f00b8ff10fe8afe3effbdff34ff84fe25fff4fe4cff74ff59ffff00;
// music[1061] = 256'ha9ff6500e701e9f3fde41ee653e7d4e499e524e673e7bde817e8c3e846e989e8;
// music[1062] = 256'h37e8bbe863e9dae874e9efea09eb25eb00eb6aeba5eb0deb06ecb2ec0bee98ee;
// music[1063] = 256'h6bebcde904e982ea08efebedb4eb82eb83ea47eec0f1c8f4ddfc1fffaefcd3fa;
// music[1064] = 256'h37f653f5bcf384f1faf96802a30342fe61f394f0dbf225f1c9f0def487fa8bfd;
// music[1065] = 256'hc401dc03a7fc9af703f860fb8afd90f4b4f09ff9d1fd1c0044021bfff6fcddfe;
// music[1066] = 256'h520c1b203f227a19891ae41e561b64153f11c40a8c060707c40a7a137218171d;
// music[1067] = 256'h2c1ec60db907510eec0a0a17732acd2c4434f934781ec90c750730071c12aa21;
// music[1068] = 256'h8d23f2174f0e1a0947079d085105f604b70a9008ef0a8d1f6e2d45243615470d;
// music[1069] = 256'h590f961a5d23c12ab33502365e2b77227919d1105616952900376d3d743fdb32;
// music[1070] = 256'h53281c30a537a836b83a0f41613c1838f5414a4d8e4c8541ea3c0e45fa45973d;
// music[1071] = 256'hf63cb844be48b64082355a2e432b4031e838f03fba40c931e931623c202ed224;
// music[1072] = 256'hc72fb439773dca36f72fb02b7d2da944b553df4dc348d84084436556a05ed156;
// music[1073] = 256'h12482a426b4aa4502e4e1a400b372545264b943d4b39603bb934b32beb2eb643;
// music[1074] = 256'h174d4d36042473258f204f1e5721aa1af41d3128e024f11d4b12630a6320ea37;
// music[1075] = 256'h5f2b95177f180f203c22651a70153721f82ab32f662ebe16ab06160e3b171926;
// music[1076] = 256'hf629a316800d4814651e361f2b0c7ef9a4f17af8a20e791264035a001602eaf5;
// music[1077] = 256'hbce10fdfe7f478ff0aee2dde34e0dfea44e956d3a0d1dae8c1ebfee405e3e4df;
// music[1078] = 256'he3e246d537c25fcde8da12d961d14bcb71d55fdcb1d6a5d9b1d882d8feeb1ef3;
// music[1079] = 256'h76e6c2e883f93d093a0fbaf83bd549cc53d53edafcddbfe85f0300174e04b4dc;
// music[1080] = 256'h62c2eec7b8e2edf7e1029b102921a70eb0d3cdb13bb68fc2ced89be12dd20ed3;
// music[1081] = 256'h05e657efade8b1e0c8ef3708d8117b1710140501eef586f9bd008d08ba0764f8;
// music[1082] = 256'h4dedc1ef65f5cc003310ba19251c14146907ab0365071707a3fe95f7fbf457f1;
// music[1083] = 256'hdaf5df0b712698367b3a392f2a18fe0bc017a524c11b8d109016021b48190125;
// music[1084] = 256'he636d03aaa35482e4f1e6112331a6d264822f611ad1360271c27ee1e7825182a;
// music[1085] = 256'hf023750b81f5bbf7ccfbf00c14269228262947221f12ae11750487ef44f4aafc;
// music[1086] = 256'h51fc8ffb88fdfb0037fe93f983f167ed92faec048b05f0fdd4f42dff7ffddde5;
// music[1087] = 256'hffd725cedfd0d2dbd3e0c6f5360653ffb3f4f3e5f2dc99e604f110edaee51ae4;
// music[1088] = 256'h2ce725ef04ec71e054e920fb60fa9fed08eb93edc5e413e7f7f7c2f84ef659f8;
// music[1089] = 256'ha5ed29ea51f4d4f51cf41afbf106b10ad807950ddd11d50f2d0e5705af00000a;
// music[1090] = 256'h6b1987227a14aa04770b6511de0b360a6a0e4f0d3209a215a0288e2780170e06;
// music[1091] = 256'hea00ca0b0617522341288c2025244529122ff63e49397c31433f47436341d83f;
// music[1092] = 256'h0938eb345835233a7f3c9736b9374f406a4a044d0443983f5e423542764bd952;
// music[1093] = 256'hc44a194b9750fe485e49e5407e1fa01d5735582eb11bdb1c5229923237354e2f;
// music[1094] = 256'h581fa2192f23ee215a1b34216c1edb0441f288fce30ae304f3f6d9f18dfe780f;
// music[1095] = 256'h3003b9efebf5c0f8c7f159f619fb8bf44dee90ef57ec0fe20edba4dfeeebaee5;
// music[1096] = 256'h94d46fd245d221d605e176dc63d05dd18ed4dbcda9cbded18cd0bcc80ec43ec5;
// music[1097] = 256'h1ec7f4c4b1c4b1c8b4c971c0a0b4efb2f1b439bcf6cd29d3bdc8d3c248ba24b7;
// music[1098] = 256'hfcc186bc98b2d6bebed04ce3a0ecb1e0bfce9dc719d416dcb4d011d124dd1ddf;
// music[1099] = 256'h87d886cf61c97ac83cd7cbedb5ea5ade9adfc0d6facf0ddd5cdfd4d51cd6edd4;
// music[1100] = 256'h64c7aabb58bebfc4d9c7ffcd2cd042d5b5e8d8f3e0edcde27edb8adc01d1fac2;
// music[1101] = 256'h5fd282e4fbe7fbec92f1caef0fe5e4e081ee4ff717f47df472f5a5e96fdbc1dc;
// music[1102] = 256'h8aec2c00f1075106680c1e0e8efc29ef6bf540fa5cff070c890bf604f208b917;
// music[1103] = 256'hc424ab1e1a1bd61a321113192628c12eff333431892f5d294b1f9e28fd330934;
// music[1104] = 256'h32395f439b42f036bf350a3cb33a8239c53c9c468f55f5591f545354c358575a;
// music[1105] = 256'hbb5e965e5f56ec54c35765585156b4533e562f57a05a95602659ad500d54ff57;
// music[1106] = 256'h2f56ec522351674b173cc42b822d4433ca2c092f4e35bf346a32ca2afd278e25;
// music[1107] = 256'h741fec1f6526702ac021ad239a286619b81d942254148416261ab71c1c1e5e16;
// music[1108] = 256'h20169b0ff20afb12cd12ff0d8f055b03950dd10bf80094fc43fe41014dfc37f4;
// music[1109] = 256'h04f5c6fb88ffc5007b00bef77ceb04eaddf08ff38deff1e98ee167d955dee8e7;
// music[1110] = 256'hc3eab9ee58eb77e112df9edb00de23e4cfda1dd597d394cc67d461dbd4d5a0d6;
// music[1111] = 256'h33dae6ded9e1e8e405f038f151f0eff524f10cee38e9aee3a9efeaf554f156ea;
// music[1112] = 256'ha5e1cde7b3ece2e44bdf2ae273f0e3f3d3e870e828e568d124c3d9c51acdbdd6;
// music[1113] = 256'hdddfcad9a7d070cdc0cbe1d053d1e6c8adc99bd7adddd5d234d00bd7afd7eed4;
// music[1114] = 256'hcdd2c0d6a7d766d423d85fd82bd4ccd102d73adde5d2c4cfb7dc51df19dc93de;
// music[1115] = 256'h23e0acdb5ad38fc986c644ce2bd7c5e25ae78de0b3dab2d3aed8bae152ddfbde;
// music[1116] = 256'h29df7cd953d9ead9aaddece21be666dc72d4c1e46be705da21dad4db42dec5e3;
// music[1117] = 256'h1ae6ace395e2b2e4fde144e5c9ea71f32310f61c6e0d3c05cd044503c5073c0e;
// music[1118] = 256'h64122214a310121712250a23f01c3c161612b21609118b11961b79221927c918;
// music[1119] = 256'h4c17091ecc07bd05af11450b9a0f3013890dfe0d3a0a9905df09850e8f127b16;
// music[1120] = 256'h5e0e4108db12d41acd184016331696147e115f12c1124012a4112214e216df10;
// music[1121] = 256'h51169e1f991bbf220426aa1a131773142319012797270e1d0e17411cdc20f21b;
// music[1122] = 256'h151bfc22282a8e26071b63167c166718d822ba2858280e2d342ae51d2b16b81a;
// music[1123] = 256'h6828822e6932e3353f2d4f2ade2dfb2cbe2f882d072471255d32f9369f36c73d;
// music[1124] = 256'h4e40b7426c46c444664848467841b543c43e213d5e42c7441e40e6318e2ef039;
// music[1125] = 256'h833f133bb93511369c34e931bd377e392824080d4911e51d4e1e4417a4129115;
// music[1126] = 256'h1b14a112f113610fdc116f123907c605ee0dcd11e616331d87133606b208f207;
// music[1127] = 256'hea025508ef0ded0815046a0fff15be09490716092502b3068b0d0a0e7c103b06;
// music[1128] = 256'hc3fb68001603cf0470019efa4bfeebfb8ff6d8f90cffed08b10b0a0026f6d5f4;
// music[1129] = 256'h89f6ddf704fc76fdfdfb47ff00ff21f8c5f648fb7df9b7f532fa91fdfafae1f4;
// music[1130] = 256'h6af1cef4e7f397eeb5ee3dfa200b2f0f680aed077306f8030f022d07af074fff;
// music[1131] = 256'h66fe0dfedefb71015f017afa6dfa95f9f3f522f54af012f5ac030f02e6f5ebe4;
// music[1132] = 256'hc6d84de011e02cd71fd8c7d897db1ddb63d6efda68ddb9d8f4d034d0ecde7fe5;
// music[1133] = 256'ha3e2c9e52ee6cfe70ceaf8e2a8dba2def6e8fee602dd7aded3ded1e12be92ae3;
// music[1134] = 256'h7ce20deae2eadeeaf5e0cbd50fdcebdf3ed801d40bd8e3df47e2cbdff7de93da;
// music[1135] = 256'h0dd75ed8dcd4e0d4a3dc80dbcad3cbd42bd560ceebd3dad8c1d2fbd84cdb02d4;
// music[1136] = 256'hb0d3f3d160d5abd518cde2cd4fd0b7d295d823db3ed90bd1c1d205e0b7e3b2e7;
// music[1137] = 256'h35f195eacbe091e2d4de34dea4e110dc83deb5e111de4fe2f8e217dc7bddc7e3;
// music[1138] = 256'h06ded9d804e36de4efddc3dbd4cd12ba41b139b2c9b482b933c0f0bce1b895bf;
// music[1139] = 256'hf0c342bc29b0f0b18fb916b95dc05dc68ebdeeb888b92fb652b5c8be3fc8ddc3;
// music[1140] = 256'hf8c286c81fc5b0c1b8bffebf94c55ec495c193c5f8c5e4c11ac621c990c34ac8;
// music[1141] = 256'hf5cdc8cd32d3e4cf2cc6afc032bed8c3d5cae5ce50d1b4cf3dce87d383d6f7cb;
// music[1142] = 256'hfdc665ce3fd389d71cdad8dc36df43d91fd230d1ecd513d7cbd403dca2e0e9db;
// music[1143] = 256'h47db31d8e8d372e2e0f4a5f507f11df3aff8e6f928f9faf946f9c7fc7dfa07f5;
// music[1144] = 256'hfbff2b0a86091f077100f7f86df99603920b7a0dff0e7710e20c8cfbe3ee63f3;
// music[1145] = 256'h96f5def4cef62bfbb9ff5cfe0aff73fff6f618f418fe80056406e70401fe6dfb;
// music[1146] = 256'h4bfffa01bc06210796090b14ca11fc08670c4911150fe80c9a0e20148b1ae319;
// music[1147] = 256'he1141f100d0e3d15c31c981cbb1b521ddc2074258124b417e21463232924691d;
// music[1148] = 256'h351f1422f023bf20e7227726ff24a62f7f33432eb730192e41324439bd311e2c;
// music[1149] = 256'h0c28ee29f735af35e7310337aa340c2dd3287c2d46414e506d4ee84a39496b47;
// music[1150] = 256'h1b4aee508f53265123505c4efa4d464f994e8f508050af4ff55349539e4b1f4b;
// music[1151] = 256'h9052d255435a1157984078374d3ddc3a2e3b313b2434c8324135a735b5397d3d;
// music[1152] = 256'h023bb133382d6133b336df328f3a953b793c5942613b9c397435a032e93b6836;
// music[1153] = 256'h46373540e43c12413540db34ea3511389f33b63586397a377a38ed3b943c393a;
// music[1154] = 256'h4c38d63552304632013732350c34e134a2378f38743ba03d43384e38f33f1047;
// music[1155] = 256'h1141b03c0a46743ce835143c0f37a13d273e82353b37be32ca325334e631d432;
// music[1156] = 256'h4631ab3aea46bf48a445ce42eb437840f33a6838d93c2946b541643cc63e113f;
// music[1157] = 256'h3f3e333c293c683972376e3a57381b37cd313f2cf6305a279012c30ff3148110;
// music[1158] = 256'h6b0c040d010d0f12c8126f09ed06b50751024efe40fb5bf830fdf30120fc72f5;
// music[1159] = 256'ha5f3a5ef61eeeaf504f720f152f2eef1cded64eaf3ea68f003e9fde168e9d8e6;
// music[1160] = 256'h1bdc93d7aed78cd4eccdd3ce37d3f6d32bcf40ca26ce14cec6c8e5c846c814c9;
// music[1161] = 256'h2ed13ecfc7c107c0ecc314c455c750c730c8ddcb6dcbb2c731c2f3c082c1cbc1;
// music[1162] = 256'he9c260c202c889c883be25bb20b941bd1cd0e1d773d386d4d9d7cddb76d72dcc;
// music[1163] = 256'hc7ccafd161d17bcacac4f8cc92d43bd327d0bbd045d47fcef5c4fcc57ad1c1d1;
// music[1164] = 256'h50cab1cc46bc02aa66accfa649a96ab15cb0eaaf03aa63a907a92aa21da2bba4;
// music[1165] = 256'h8ca3409f83a1c3a08b9b889f399dcb9e3ba667a2189e58a041ab46abab9c329d;
// music[1166] = 256'h03a5eda62aa420a0e39c9e9bdc9e039e5da18ba8cea5f0a356a296a5ffaa25a5;
// music[1167] = 256'hffa334a4a29d2c9eada3d7a5d5a1699da1a2fcadd2ae56a9deae87afa8ab1eb1;
// music[1168] = 256'h90afa2afe7b3deb05eb69db68fb1f8b98cb680b103b87fb3bbb3beb750b86bc8;
// music[1169] = 256'head3c4d119d180d14bd637d931d908dadbd5d9d4f0d68dd46cd50ddcfbdfacdf;
// music[1170] = 256'hdde0e0df6dde84df48e2caeae6ea7fe85aea28dab9cf01d14ccb5bd303d9ebd2;
// music[1171] = 256'h82d3a1d2f7d4c8d9f4da2edc74d9a7d7d2d506d4c1d7fadadad785d72ce17ae4;
// music[1172] = 256'h03e3eee54fe277e28fe6d2e37be47dedc5f08de8cde824ee2aef3ff06ae857e9;
// music[1173] = 256'hd1ef3aed2df26ff379f39ff653f4c9fa2efc04f8cafdfefb14f42bf2fcf2bbf8;
// music[1174] = 256'h2303a5053f02170114008e05070c1e09f006b70d3115420f1b0b2514e819ac1a;
// music[1175] = 256'h9e19e716c2197a20941fd121cb33b03c093f3842a83d9d431d474740c241ef41;
// music[1176] = 256'ha2439747934a1c54f15bd75bb05c695f035b575f126d8f6b3168c4661b635e5e;
// music[1177] = 256'h61523552db54a44f5751a64e7e4fb354bb51aa572e5df155d7505451f355065b;
// music[1178] = 256'h785c0a5d835aae56b957045b055e245f9d5bc058a05d20627a5a7256dd613f67;
// music[1179] = 256'h8a618c5efc5d275f8d61ca60a06129616959185aef5f9a5be3574b59a85d2d5f;
// music[1180] = 256'h905e0c61af57de53a158b551ea557e58465364595b535b4fae561958925b9256;
// music[1181] = 256'h6d4ed4501054ea54a552f355655a5356d44c1242da41863f883e5652b75ee65d;
// music[1182] = 256'h3e5d4c58c257f9577e541c52355265545d54ea587d5b0b53ec51415a915e885c;
// music[1183] = 256'h135abd5833557c52954f4c4e99487e37b7329539a6353b2fac2d573108364b2f;
// music[1184] = 256'h32262927e829332b512b3c288d28e9279120721df7215b28c826191fc91d061f;
// music[1185] = 256'h19201121a31e561c6d18cb17bf1cbb1a1f18381de917090fd2155b16e30fd813;
// music[1186] = 256'h22149715df17a30de107f20aa50d3710550faa0b4808ac038100c5075f0e1309;
// music[1187] = 256'h5e0784071d0266038306e002a6ff47fc33fb66ff53ff1901ce042a036c0160f5;
// music[1188] = 256'h9aeec7f7c1f3e0f36e066410c60dc408b4064204e300b2fe05000103c4ff47fe;
// music[1189] = 256'h8afc70fb8500cdfa0bf74cfb75f9ecf4dcf0d6f4d0f49dec88ed17e841d61dcc;
// music[1190] = 256'h33d2ced2bac803c964cb7ecf47d10bc612c2aebf5bbb44bbf6b82dba3bb70eb4;
// music[1191] = 256'h61b7a3b541b512b695b308b107adbea9bbab87b389b43fae47ada0adc6b039b7;
// music[1192] = 256'h77b193a4b8a1f3a51ca765a48da4a8a59ba3aca78ba7579fdf9f469cf098a7a2;
// music[1193] = 256'hada35da048a2ce9f399eefa06d9e0999969b4b9f5fa0c2a1e59d789c9e9bfa97;
// music[1194] = 256'h289c9f9fa39a49964e9ab49f339a5694d19467948f9bedada0b590aedeacf8af;
// music[1195] = 256'hdcafd0ac09a908aa7dab0cac8ca9b4a591ace0b141af43ac2ea951ad55afeea9;
// music[1196] = 256'h01a864aa04b29bb026a3c89b0c961c91e4915893bd96a1963d92d9929b958896;
// music[1197] = 256'hc1977d976e92408bab8c0096c59698921c93d08e048c8c8f2d8fee93999e3aa1;
// music[1198] = 256'hb49cd99cb5a3b1a25da17ca71ba2769d97a2869f8a9e79a32da160a0e7a5e7a6;
// music[1199] = 256'h60a2d8a091a2ada4e5a5dba3b4a693acf7a6b1a24ba9ada9eea5d6aa00b164ae;
// music[1200] = 256'h01aa82ae7bb14bab73a9c0ac1eae12b0c5b051b163b4a6b479b187afd9b31eba;
// music[1201] = 256'h9fbbaec5dcd2f0ceaacc9dd3b6d08bcc0dd32fdc87dd0bd838d70cdb5cdbe1d7;
// music[1202] = 256'h1cd77fdd2bdf26db63e3a9ea18e527e605eab7eccbeda6ddb5d02cd161d095d7;
// music[1203] = 256'h46daf5d62be002dc13c9d9c8c7d075cf1ccd6fcc66ce0ed525da30daeed52ad5;
// music[1204] = 256'h89d93ed64cd481de67e2a4e0a4e661e8f9e53be9f1e7abe7c0ed7fecaaeb99f2;
// music[1205] = 256'hf3f4d4f13af351f7bdf5e9f459f7b0f58ef048f392ff0a0010fe4e0733043afe;
// music[1206] = 256'h84ff5fff74061109f406150c750a07061b0be50e950ced0aa50bfa0f4213e011;
// music[1207] = 256'ha913041477148317bb133d16fe190313451d9d33c738f7366d395b3af6390837;
// music[1208] = 256'hf136fd3d853ee53b803ebc3f8a43004623451845a9408c3f6043fc47a44d2a4a;
// music[1209] = 256'h7b474c4ad13da82c5c2cc833ad384038bf33d635d93a0c379c325935be387939;
// music[1210] = 256'h813b433ec53d793cd23bbc39d039f23cbf3bd6367f39ff3fa03d293de642d33d;
// music[1211] = 256'h203b67438e42f03fa84495478e441940f3459146423e5a4252459245cb4b8b49;
// music[1212] = 256'hd147534c494afe47c64a014aa249424eed4f434edb4a5e4784466548eb4f1052;
// music[1213] = 256'h4e4b8c49604bf34ad54be1514c537c4ef0517f54844c4648f64f4553ef4c2059;
// music[1214] = 256'hc96c176baf67156bd168d8682f7073702e6977676f64f062306bf46dbb676565;
// music[1215] = 256'h886a8f6d68682a679370ea7349682963f7633a57cd4d9c5062515f517a51974f;
// music[1216] = 256'hdb4db14b5c48ca467449ff4c0c4efb4bf74b264fc04abd450f49b349c8482149;
// music[1217] = 256'h6c45ac3e143a3a40734520423f45a6455342e0456a422a3e7041e840473dbc39;
// music[1218] = 256'h3e3b263f4b3a103768398635e034823b66380c325a350f384a349c31f8332d34;
// music[1219] = 256'h4030d42ee62bcf276c28e927aa25ea2aff310e30682f5933d02fc52ade2a3e2c;
// music[1220] = 256'h042f3c30552c56286024732303353946ec3e0239ee39e834bd36163afc38bc39;
// music[1221] = 256'h5536d834c138bb35a02faf2f4a31fe2fe030cb329a2d882dc931d127ad22dc25;
// music[1222] = 256'h52194b0d6d0f740fdb08f3053d080f0a32098b032f03790879035afc62ffd504;
// music[1223] = 256'hb7ff74f937fe26fe62fb3afae2f4aff4bff288ef76f19fedc2eacfefcaf3e1f1;
// music[1224] = 256'h1eefe1ebebe95ced8aec76e878e450e361eb09e942e34de91de9cbe53ce2bddb;
// music[1225] = 256'hbddae2d7b1d467d5f7d3e4d466d5face27cd18d213d434d294cd77cbfecb05ca;
// music[1226] = 256'h2ec928c7c6c71ecdc0cc2bc9dac50ac582c1ddb94cc0a8c56bc3c7d2e3dea0da;
// music[1227] = 256'h3edc16dd3ad685d59cd830d5d7d1c3d168d1ccd5c7d81ed522d303d303d434d4;
// music[1228] = 256'h61cffacac1cd3dd2f1ceb1cda6cc88bc79b1bdb3e8b3fdb275af30ae98b172ad;
// music[1229] = 256'h03ab8eb103b1e5a99aaaa6ab99a751a72fa926aacea9d5a84ba73ba3d2a26ba3;
// music[1230] = 256'h5ca376a3819e299da29f2ca14ba4bca57ba5a09fa29b819e069dc7a02ba8dba4;
// music[1231] = 256'hc59ebc994996cc9b9ea1e19a4c96a99ca79e5f9d309d5a9c019c969817944893;
// music[1232] = 256'h74969999aa9bce9c6398669a65a2769f199c389ed79b7899bb997e98df984399;
// music[1233] = 256'hd994929239922497f8a97db731b6aeb3bbb1acb1e6b1b9afeab1f3b32bb25bb7;
// music[1234] = 256'h71bc4cb7b2b434b673b75bbbf7bb17ba83b83eb95bbc95bed2c9e3c879acce9e;
// music[1235] = 256'hc3a343a352a4f9a8a7ae38b1b5b2ddb63db317afb1b048aeefac43b0c0b3cab5;
// music[1236] = 256'h3bb459b0e5afd1b491b7a6b462b279b3efb303b33cb619ba37b80eb8debbb4bd;
// music[1237] = 256'h9abdacbadfb6b9b895ba00b92dbd32c249c05abf76c150c442c6b3c362c3dec8;
// music[1238] = 256'he2c9cfc48fc387c896cbf2cb15cde3c8fec5a6cbabca07c58cc801d208d4c3ce;
// music[1239] = 256'he2d327d688d180d8aed7c9d765dd13d71edb64d91fd7cdef9cf81ef757fdf9f9;
// music[1240] = 256'h4cfc1efc8af5fff9adfbecf635f9cafff60083016b05480619077e0733025cfe;
// music[1241] = 256'h2f000603510f481dd5111a004efedbfefa03c90bc3082e03e3067d099008660a;
// music[1242] = 256'h710482029c08b405490ab310620c9c0b4d0b5c0b610caf0aba0ab80c59118212;
// music[1243] = 256'hfe0ef9091e097714cc19de12ab127316ea148c114415041cdf18d116601d7a1c;
// music[1244] = 256'hed18e71b9c1b481b091fdf20ef1fa81ff1221f221c222327cd233a23b625951e;
// music[1245] = 256'h511f382551226b23d4292627d421f224dd27f72aed2b9c2476247629bd2bff2e;
// music[1246] = 256'h232cfb2e6a40ba4c414c13472a447b4626482941e63b8542d144de407140493e;
// music[1247] = 256'h1c41404824472845c4462547fc47d7485e473349b74e1545d72f472c2332fc2d;
// music[1248] = 256'h9730953809350e36ff39b933a933b4337a328a3aa037cd34393b5b337c2e6b35;
// music[1249] = 256'h5e346d32b636da39a23ac438df32ec305d34b435cb348f34a138173857301d32;
// music[1250] = 256'hfd354e353837463720373637a8335f3295389d3cbe3741392c3c27366935b738;
// music[1251] = 256'hb839e23a213cff3b6e36e832a2342e35f335ec343a32b5327031d02f7c33c431;
// music[1252] = 256'hab2df7305a319a33f1369f33d732582c782e84465850934ba74c5b4aa045c144;
// music[1253] = 256'h1944d74297420f4367463e463642a746034922452447b746a241a73f9a402d40;
// music[1254] = 256'hf9412644f13463217c1f2826ef2a66287828902df12734219d232526ab24d622;
// music[1255] = 256'h5f2373238a2377210d1de21c851c201b841d7d1f281fb61ec71fc720af1db81b;
// music[1256] = 256'he51d891c431c2120de1d641a3d19211642165c195d1b4b1b061c291ecf1ba718;
// music[1257] = 256'hd518271cbe1cce175919531ac713e6147b1a5c1a541607153a174214f60f7915;
// music[1258] = 256'ha61b91172217aa1a8a1798181e15820ea215eb1760143b1373113615ca12ad12;
// music[1259] = 256'hf722242b5828df27ac260227aa2a5c2b3729ee256421af217124af2331253629;
// music[1260] = 256'hec2ab828812508246f23b42391219a221225b7165d0604053704e404a10ba50c;
// music[1261] = 256'hbe070e051b04a20257045f073e05b5013e004500000279ffbbfd8302c70090fa;
// music[1262] = 256'h4bfa86faa8fa05fd20fe30fd83fd48fcf0f63ef6ccf853f9e6feed04f9032c03;
// music[1263] = 256'h32052d047a00adfe8400ec04f605d40112fe0dfd19fd71fbf6fa33fe3b012202;
// music[1264] = 256'he6ff39fceff88ef5e7f32ff42cf77ef9faf683f519f7e1f74df66af58ff783f7;
// music[1265] = 256'h8bf6def67af4fbf4acf560f014f53803f1067b05c306fb051006cc084f090106;
// music[1266] = 256'h04041304bdff31fe27053907b603f1039c049703f1ff02ff9e04200105fdaa00;
// music[1267] = 256'h63f303e3c0e31ae70ee9e1e68de4e4e62be53de554e564e146e40ce84ce6afe4;
// music[1268] = 256'h15e125df1be0cbd647cb43cc34cea9cd05cfaccfc6d004d0dacda0cd4dceeecf;
// music[1269] = 256'hddcfe5cc24cb1bcec2cf6ccc2fcc40cd9fcb57cb20cb53cbcecb7dccb9d143d2;
// music[1270] = 256'hb2cab8cb8fceb6caa2cea0d126d074d366d05ecc32cdadcd32d118d01fcd45ce;
// music[1271] = 256'h94cd18cfa7d17fd1b3d1b3d1b3d0ccd0f9d2b3d315d6d9d679d3b8dd6eec95ec;
// music[1272] = 256'h92ed7bf198efb5f07af3aaf0d3ec21eab8e91eee4bf269f35ff3c4f2d5f2eff2;
// music[1273] = 256'he8f2eff373f631f69af02cf1a8f5efeb92dc9dd723da0adee2dc0ddb16e11ae3;
// music[1274] = 256'h03df83e07fe1c0dfd2e0cdde55da57daf0db52dc75dcd6da62daf9dc97ddd9dc;
// music[1275] = 256'h2edd78dda5de57de89db20de6be31dde72d7cfd9dbdb00df10e143db4fd961dc;
// music[1276] = 256'h6fdcf9dcc1dec1dcbed8add854dc08deb2da7ed913dd47deabdee4dc6ed81ed7;
// music[1277] = 256'h99d53bd58dd854da12da26d945d642d53eda61dc04d94cd66cd6f5da55da3ad7;
// music[1278] = 256'h82dad7db7dd9ffd5eadc87ec57eea7eb16efb9f182f071ed21ef26f06bef04ef;
// music[1279] = 256'h74eb27ec77ee83ef81ef0bedd1f012f413f09bf02cf266ef18f2d8f021e0aed6;
// music[1280] = 256'hb3dbb1ddead8c8d4fad7bcd952d76bd844d8e6d981da40d674d8dfdb34db31db;
// music[1281] = 256'h18d897d581d7f0d54cd3ffd364d291d1b6d262d409d85bd9e0dc5ede37da3ddb;
// music[1282] = 256'h37d9d4d5bada16ddfada92d826d850d8f6d70dd86ad2c4cff3d6a3d9b5d5ead3;
// music[1283] = 256'h18d7f0d9b3d6ccd169d41bd94cd593d326d530d10ed1fdd121d1e2d2b5d0eed0;
// music[1284] = 256'h1ad5ddd3ead0a8cf3ed1c7d46cd7b4dc3ae266defbda07ea2bf994f8ebf896f9;
// music[1285] = 256'h8ef6a0f86bfc3efbf9f6d9f877fb89f954fcecfb73f9a1fe15fe61f817fd1505;
// music[1286] = 256'h800204ffb7006701e4fff1f148e77fed39ea6ce5bce982e97ceb99ec3eeb52ed;
// music[1287] = 256'h0eefc4ef49eec1f00bf490ed5fe8ebe9d2ecedef67f1ebef00eee5ee28f178f3;
// music[1288] = 256'h71f3b5f1ecf3f5f59ff5e0f4a2f48ff82ff6daed61f237f741f2aff5d9f9f0f4;
// music[1289] = 256'h86f4d3f7c5f8d2f7f8f6c9f741f64af6cef9e6fa27fb82fcbcfc83f7d9ef5bec;
// music[1290] = 256'h3aecb3eee0ee22ee78f2d3f45bf39ff11bf1e4f379f4e1f2eaf4d3f67cf602f7;
// music[1291] = 256'hacf4f9f41503d30f090fab0e3512b912e011041385132a12e712e413cf12a613;
// music[1292] = 256'h58152214a013f617ad1c911d731aa617261d75238b21ad1a260d2506b70c460b;
// music[1293] = 256'h1809c40dc1084b066b093d08dd0bf70e4f0e1c0e050c3d0e8c100e0da309b508;
// music[1294] = 256'he80a250d760fcc12c3126911a50f1c0fbd12d5154a17041743148a120913bb14;
// music[1295] = 256'h0a139c103713a61506197f1b8019c419c81633144118d718631ac2191415041a;
// music[1296] = 256'h221c86173a195a1b621a441a481bc2195717181da7239623b523cc21b21e8d20;
// music[1297] = 256'h9721c320d2208222012551230d224f206d216d32b93d783aee3b403dec3ce73f;
// music[1298] = 256'h1142d440283db23d7d3e5c3d393f753ed93c92408743c7414e42be438f43f745;
// music[1299] = 256'h2e459646b64516344d2b962e182bf72bd72ea02d6c2ca62a672b4b2cd82eb431;
// music[1300] = 256'h9c2f98306732b7309030bc2eef2dd93002312a309330e12f802f88314333d130;
// music[1301] = 256'h8a300036d3371135d1345c351833a930ca2e8f2e6d3114315e2e762d072fc933;
// music[1302] = 256'h6733a9304732c7305a2d4b2df4324534042fb332f3330d31043448319c313735;
// music[1303] = 256'h6a33a8346133b33379377133e130d130922eac30a831132ffc31f3342030e431;
// music[1304] = 256'h613fb445dd4379471b4b7d4a5f4c524cd2489248b5481847ca455b44e343dd44;
// music[1305] = 256'h9a44b5453d4b6b4df44b4f4c404aea49424c1546e138e53109344133092ffc2d;
// music[1306] = 256'he02c4c32523baa3bc83a913adf39c53dfa3d183a5e3a913b8c3bee391c371937;
// music[1307] = 256'h6c371037d13690339c33563861371d345a345a3415344f328230203443378434;
// music[1308] = 256'hd5317331be2e642cfa2d1c2fdd2ff62ed52c292e1f2c172bd12ea12b9d275726;
// music[1309] = 256'h612401262827f2275828e1267b27ba2718277025e622b1231f25e0233323c525;
// music[1310] = 256'h7d247b1f2f1f092283246220061e6c2aeb341a3758382037d534a53104312f31;
// music[1311] = 256'hb92f0c3152318f31fe300b2ca32a672af322a31a801a3d1c4b1d3c1e911b3f1f;
// music[1312] = 256'h961b5307b7016a04df006701e20098011903e7ff90fd14fcf7fb74fb38fdb001;
// music[1313] = 256'hd2ff77feb7fd33f970faa8fb82f9e3fb21fbf9f507f40bf2b0f1e0f4f9f4d5f2;
// music[1314] = 256'hd7f241f46ff223f065f14ff1baf24ff262eba0e93dea06eaa5eb98e98be88ae8;
// music[1315] = 256'hece590e620e8d8e494e0ece233e5c9e1e1e0bae19ce3b4e66ee310e05de1a1e0;
// music[1316] = 256'h35e04fdf90dc0fde76dcd6d8eddbc1db4ed951d965d844d88ad51edb96eb84f1;
// music[1317] = 256'h90ee5fec0cedbcf00af0a1edefece8eadcea81ebe0e790e613ebc8ec21ecd8e9;
// music[1318] = 256'hb7e52ae577e45be693e98ae802eba2e396d2a5cea4ce30cdcbcef1ccbdcb49cd;
// music[1319] = 256'h3acef0cc36c9cbc6bfc6edc856cac5cab7cc86cbb6c87dc810cacfcad4c7b8c8;
// music[1320] = 256'h87cb82c606c487c619c5f6c386c31ac2e4c3bcc5b2c58dc6c6c5edc3b6c3d6c1;
// music[1321] = 256'h25bf86bf6dc0b8c01cc159c0f7c00dc24fc08abeb4bdfdbef3be18bc18c0d7c4;
// music[1322] = 256'hbbc25abf54bdabc01bc2b0bf7bc0c9bec1bdbdbdedbcadbeb2bdbebdd5bdc0bc;
// music[1323] = 256'ha8be6bbe9fbda7baf2c0f2d2fed638d540d77bd5e5d574d56dd558d80dd9b3d7;
// music[1324] = 256'h45d6c0d654d868d954d775d5a2d5f0d413d835d55dd18dd6aad7f9dbe1d7b4c5;
// music[1325] = 256'h71c374c4b4c124c568c318c2c5c127c0d4c151c0e1beabbf04c029c233c2f6c1;
// music[1326] = 256'haec4bbc5f6c487c40ac5c5c6aac688c44cc330c430c5cdc546cb5acf7ecc9fcc;
// music[1327] = 256'h5ccc89c913ca8ecacbccc3ce4bce40cf50cf49d112d213d403e2ceeab0e6e9e5;
// music[1328] = 256'h51e66be5d1e860e9c4e60ae881e8eae7b6e861e86de85be648e3d7e25de33ce4;
// music[1329] = 256'h24e1bbdf29e3e4e11de10ee1cbddbddbdbda7cda88d761de7df017f482f16bf3;
// music[1330] = 256'hd4f04df0a9f0c6eeffeea0eecbec80eb22ec67ed92eebdef8af0e5efc3edcced;
// music[1331] = 256'h7bee25f0ecef1fee8ef186e931dcb4dd24ddd4dc5fe0fedd03de0dde14de8ae0;
// music[1332] = 256'h73dff1de4bdf07e0dbe067e068e02de14be45ae5b4e374e6dee8efe578e257e1;
// music[1333] = 256'hc4e2efe5e7e007d75ad7fdd957d9e9d904d95fda8ddddfde07df30dea3de43df;
// music[1334] = 256'h3bdf73df63e14ce325e09edecbe0ffe195e5a7e745e69ce6c2e51de5a0e8d5e9;
// music[1335] = 256'h35e88ce928ec12ed01ed22ee4aee16edfaee1cef23ef4ef231f203f2f7f059f0;
// music[1336] = 256'hc8f3a1f3befbba0c0c11640e0010c112f413831433163f16271504152b158515;
// music[1337] = 256'h9517d61ad31a701aac1a4e19c9191219a0187b19e519a71c2015e408f708ec08;
// music[1338] = 256'h4005ef04e5075e0bc009e809630b4809dc0afc0cbf0b9f0b3d0e27119f118c11;
// music[1339] = 256'hc0118e134a157914c614b512990e9f0fd811d4103e10b7114c123413a4157216;
// music[1340] = 256'h55163616e5166218fb19471bb618ce15b6164b171216a21491145615e216f717;
// music[1341] = 256'hba182b1b8d1a7818ab19c21a311b341b041bb319171a7b1db91c2d1ba51b961a;
// music[1342] = 256'h921a1f1b161b781af21a911bd31a59197316961f4f307c3351333935d4348536;
// music[1343] = 256'h69354034483730381d36bb35ef36993673365636df366d388b361f35bf354336;
// music[1344] = 256'h8e366d370d37b52a0220cb240b25c5227225db23172333233b220b2446252421;
// music[1345] = 256'h411a481bd91f3a22a1274c29c02adb2e082d472b7229ca25272494201a1ef31c;
// music[1346] = 256'h2d1aa2199a192c18f218e71a0b1a541ae51cf61c891d211fc41fff1ff41df41c;
// music[1347] = 256'h1a2034236e224a21142232226c2324253225e22521271a2870281e29502ac42b;
// music[1348] = 256'h3a2d152e3330363103310a324131e5306b311231f530423121332c35a1332831;
// music[1349] = 256'h023c4a4de54d4c4bd84b4f485e4f4f586b576e562255d9539c532453ca52f151;
// music[1350] = 256'h23529e516a4f534e3a4efc4def4c5f4b734cc04a133dbf31fd322033a7308f2f;
// music[1351] = 256'hf22e5d2fc02d062c5c2b54290727092682268e247122e6247627ca275327b526;
// music[1352] = 256'h4d263a25d7232622a91f351ef31d0d1c501a371a5d198a180d18db173318ea16;
// music[1353] = 256'hd015ea15991560156b13c80ece0b210b570a930a810a54092c0982087708c308;
// music[1354] = 256'hc907fb07b007010693036101c2011901d3ff89ff2efe66ffedfdc7f229eb84ec;
// music[1355] = 256'h60eb27eabaeb4aeacceab6e910e7fcf2ce002c01cd00cc01d200540168013901;
// music[1356] = 256'hfd009cff23ff17ff18ffb1fe70fd1afeb4fe86fe9fffb5feaffee1ff4efe5600;
// music[1357] = 256'h16fe12f0ade826e9c2e7cbe9d0ea65e8d3e803e95ce843e898e7ffe6cbe6c0e7;
// music[1358] = 256'hc7e764e813ecbced6eedbeec92ec24efc3ef38eec0edcbeb69e94be943e985e7;
// music[1359] = 256'hf7e651e84ee8b5e723e887e8e1e8f3e9f1ea77ebfeeb8cea96e712e75be8ece8;
// music[1360] = 256'h36e9e3e968ea6cea1aea67eaa0ea30ea72ea3beabae9d3e9cae888e81ce90fe9;
// music[1361] = 256'ha5e978e900e9bbe99de9e5e9faeaf9e9d3e974eaf7e88ceaa1e99ce81df77e04;
// music[1362] = 256'h4c0432043004d903c004bb045f05510545056e05e604c104380444049d04a104;
// music[1363] = 256'hd1042005dd04b004db04b1030f06c70397f35deb02ef21eec6ec58ed79ed95ed;
// music[1364] = 256'h77ed4dee68eefaee68f0c9efb2ef3af102f268f21ef36ef3d5f3a8f384f278f2;
// music[1365] = 256'he0f26df2c8f1c6f0fbef85f0b4f092ee0cedaaeda2ee18ef3aefb4efffefabf0;
// music[1366] = 256'ha0f0c2eea7eef0ed19ec80ecd0ec61ed26eee6edbfedb6ed03ee36ed3cedebed;
// music[1367] = 256'hdfecdeed9cee31ed27ed52ec20ebebeb05ec75eb25ec6febc3eacbebbfea17eb;
// music[1368] = 256'h75ebb8e9e6eb55eac5e9def75f03fd026a028103f303390317039b03f3027303;
// music[1369] = 256'h6d03a5026c03b0020d02a502c9017102af03f8020f04430477022805d30101f2;
// music[1370] = 256'hb2ea47eed4ed47ec9fecdeec93ed17eeb9ed9bec8bedf7ee1df0b2f3acf3b4f0;
// music[1371] = 256'hbbf57100db04aa02f101aa02ac02f002a602d7011e011b00bdff6e013e021700;
// music[1372] = 256'h8bfe9cfedcfe50ff6b00ea00cbff55ff040076009fff15ff0b00bdff6fffc2ff;
// music[1373] = 256'hc3ff3f0055002e01a10054ffd9fff2fecefe6fff87feb3fec4fedbfd77fd8ffd;
// music[1374] = 256'hd3fc22fdaffd83fc81fcebfb14fceafc0afc89fd16fbb6fc260c7c15bb14cf14;
// music[1375] = 256'h2e15ec1446147f145814f8134e14d513bd1370140014d6120f13e612c512a013;
// music[1376] = 256'h3f12a3129d11900dff0e230b13fc97eee1e7c1e7dbe803e72fe6b6e739e9ece9;
// music[1377] = 256'ha2e958e9ddeaeeeb5bebdbea15eb8fec5eed3fed10edf8ecb1ed79edbced2bee;
// music[1378] = 256'h8ced08eee5ec69eb24ecd3ecb5edbbec70eabdea00ecc4eb11eb52eb2fecf6ec;
// music[1379] = 256'h6bec9ceaf9e95aead9ea12ebc4eaabea06ea53e9ffe926ea27ea6decffede6ec;
// music[1380] = 256'hbcebb6eadfe9ace9a4e9f3e90de9c2e71ae882e7ebe6e0e7aae712e80fe844e7;
// music[1381] = 256'h77e81ae6d9e82af80901f6ffa9ff44006100a5ffffffb4ff41ffb1000800f9ff;
// music[1382] = 256'hf400dcffafff810018012b01c300fbffa700a6007dfff10169fb20ebd4e56ce7;
// music[1383] = 256'h0de885e9dee826e790e668e7bee787e7ace85be99ee900e92fe8bde8f8e9ceea;
// music[1384] = 256'h83eaafea6deaafe9eee9dbe918eaa9e984e9c2e90de889e701e8bee8bce9e3e8;
// music[1385] = 256'h34e8ede691e448e366e3f1e51be805e715e6dfe6fde624e7fce7a3e852e9e9e8;
// music[1386] = 256'h6be842e8b6e7e4e708e7e6e6bbe7cde660e619e6b6e578e5f7e42de552e40de4;
// music[1387] = 256'h3fe4efe3f0e31ce329e456e4c8e35ee5bae248e76af76cfe0afd03feb4fe70fe;
// music[1388] = 256'h9ffeeefee3fe7cff9200270085ffc4ff9aff56ff32ff60fe03feb5fdaafc7ffd;
// music[1389] = 256'h1afd64fc38ff10f706e7afe4c3e618e677e82ce566e17ae471e573e733ed77ee;
// music[1390] = 256'h52ed3aee7aed1cecf1ec0ced2dec6deb71ea07eac0e9b3e9abe976e973e944e9;
// music[1391] = 256'h30eae4ea19ea66ea45eb88ec17eeeceb26e997ede4f350f457f3d8f2bcf006f0;
// music[1392] = 256'h70f064f05ef172f29ff3aff5c3f668f80dfbf1fbadff6509f011a313c312cb13;
// music[1393] = 256'hb313a7128b126012c912a312501208123d1120112c10dd0ff10eba0d820ebe0b;
// music[1394] = 256'h33106d1fe82442227b22f2221622ee200221cb204820d4205d20891fe21f2b1f;
// music[1395] = 256'h981daf1df41c1e1c971cdf1abf1b7c1c1b1b591d801457042c02c8039401ff01;
// music[1396] = 256'h0303bb02bc02e8037204d5046905c00478042104cd042e071b085408af085108;
// music[1397] = 256'h90075a076f074507de0774083f08e70753084c091208ac069506080677066707;
// music[1398] = 256'h6f07f60236f9c2f4f4f530f452f366f518f555f48ef453f490f546f6c1f5e0f5;
// music[1399] = 256'h25f5dcf422f525f52cf56ef490f47af4eaf353f459f481f5e2f6baf6f3f665f7;
// music[1400] = 256'hdff6a5f6e7f757f7f9f701faeff732ff0410bc15ff13c11462155c152b167a16;
// music[1401] = 256'h4f1684173d1865198e1b361b5c1ae3196819fc184e18871741162317b3168f16;
// music[1402] = 256'h7f191e0f5fff93fe5e00edfe470071007d01b704fc032b02920286022b04c604;
// music[1403] = 256'h5003b705180742060e07130785070908c50715088f07bd0746093e0a410af509;
// music[1404] = 256'h550ad70ab7080a065e07f9088e09f10a0d0a980ae40bb0098609f50a0f0b3e0b;
// music[1405] = 256'hcf0ad00a360b370bc80b150c540bda0aa60afc09740a3e0b210bd50a260ad509;
// music[1406] = 256'h5d096609160abf091b0ab8094809d30983086707b305bc057f07b005070ec81e;
// music[1407] = 256'hec224421e72240224721f8210f22582243235d2359238123dd231d24d1232e24;
// music[1408] = 256'h65232823c023c62252241b24b92305250819a00bf60b850c510b560ca30c6d0e;
// music[1409] = 256'hbf10e80fdd0e360f9b0d940d4c0f231068120913e51275151217e5118909c50b;
// music[1410] = 256'h4c11eb11ed15ba18b1192e1bc2199d1927184f1428124c108b0f0110470fbc0d;
// music[1411] = 256'h810ce10ab60aff0bd50baf0c6e0db50d8f0fff0fba107411d610c5126b17f819;
// music[1412] = 256'h3518e217a018bd1735195a1acc1a7d1c431ef91f8221c7230c250827bb29922a;
// music[1413] = 256'h3e2d142ee92e9f305f2f1039bf48ad4beb49c24a634a5f49e74855482e49b54a;
// music[1414] = 256'he349da47ec463846444366450f4f76522552c452ed50af515650d04f4a500142;
// music[1415] = 256'h413423349b33e6322234f9331a33f93095304b31492f9a2c8a2a192a6b2cdb2d;
// music[1416] = 256'h982bd6284d27b824ed2221220f20291fc21e7a1d171d981c521c731ceb1ade18;
// music[1417] = 256'he8185d190f188517b2173a17df160e1477105510d910df0fbb0e1f0d520bb40a;
// music[1418] = 256'h9f097607160675041103c8026c012f00bdff51fe22fdeafb40fa88f945f83af7;
// music[1419] = 256'h5ff7def667f65bf52cf4cbf337f30ef3a0f177f02ef072ee6df1ccf634f65cf3;
// music[1420] = 256'h3af2cff1e9f04bf04cf0cbef0eef96ee7ceed8ed76ed85ede5ecb2ecefeb03ec;
// music[1421] = 256'h89ebd0e98cea37e934ea33eabfda1dcf00d14cd079d010d328d276d12ad142d0;
// music[1422] = 256'h59d1d9d2c8d11bd1ced2b4d485d5f3d448d452d4aed5add775d7c1d65dd66bd5;
// music[1423] = 256'h65d50fd5c0d46dd48ed2fad1cfd2b4d233d3a1d494d47cd35fd303d302d244d1;
// music[1424] = 256'h03d1b3d116d2d5d1c2d1e0d126d2d0d1a1d1b7d12dd12dd175d1ebd145d25fd1;
// music[1425] = 256'hfed0c1d0edcf34d0d3cf37cff2cf74cf4dcfddcf39cfe6cffdcf10d04bd199cf;
// music[1426] = 256'h76d001d1a8cf0ddc09eaebe93fe98deadae995ea1aeb1cebb1ebe7ebc5ebb8eb;
// music[1427] = 256'h65eb7aeb1ceb3dea94eae4e95ce9c4e97be95cea81e9a6eaa5e993da3cd051d2;
// music[1428] = 256'ha3d1d2d121d3dfd1f8d1e7d1c4d1e6d145d203d5a2d778d71bd796d80ad91ad8;
// music[1429] = 256'h56d85bd843d820d99ed888d735d8c6d82dd97bd951d718d6d2d78ad8e7d8dbd9;
// music[1430] = 256'h10dae5da18db0bd8cfd504d72ad72ad6dad628d792d670d68dd6dcd6d5d65cd6;
// music[1431] = 256'h5fd6a3d6cfd615d716d726d76ad774d7a0d7bed7e6d7bad7c0d7b1d895d8a9d8;
// music[1432] = 256'h5fd8e2d627d87ed81dd8dcd904d9aed9fdd915da39e71ef477f356f374f597f4;
// music[1433] = 256'hbcf4b3f5cbf51cf659f659f6a7f6c0f6d5f6e6f664f723f8bbf78cf80ff9c1f8;
// music[1434] = 256'hf7f965f91cfb02f9b1e9b9e0bae3b8e4b3e4a7e4cce391e368e369e35ce304e4;
// music[1435] = 256'h98e5dde709e9c7e878eabaeb00ebf8ea72eb96eb2bece4ecd3ec35ee5cee3cee;
// music[1436] = 256'h24f6ecfcacfcdbfd98002303ab03dc03e504d602a40196006bffba0183019900;
// music[1437] = 256'h7201c1002401a6016a01e001fd011c02ff0111021502ea011a026c0144019e01;
// music[1438] = 256'h5c0127020102ff003901e2003001d70179011a02bd01ad01b0023302b6031303;
// music[1439] = 256'h9403c8118b1d0c1c2f1c211e0e1d021d4c1d4b1df51d271e401eb11ebc1edf1e;
// music[1440] = 256'hc51eeb1e541fb51ef01ec91e971e2c1f751e18215d1d0f0de306eb0a5a0ac309;
// music[1441] = 256'he2093409c6096a09b6087c0ae50849ff5efac9fd28ff57fe38fdbefca1fcd0fb;
// music[1442] = 256'hf2fc0dfd96fca3fd3efd8dfd7efd08fca6fca3fd2dfe23ff73ffd2ff4200a8fe;
// music[1443] = 256'hdffc27feedfe3cfdf5fce8fd9efd3cfd37fdd4fcd1fc0dfd1ffdf8fc8dfc1efd;
// music[1444] = 256'hfffcbffcd8fee8ff49ffb1fe06fe4bfe2bfe8efd90fd61fd21fd93fd3bfd60fc;
// music[1445] = 256'h27fd8dfc0cfcbafd1dfd92fde2fc7efec40d2d18ed15dc169c17881648170017;
// music[1446] = 256'hff168e17fc173c185d186c183d1844181718181857188f186718f718cf196018;
// music[1447] = 256'h631acf157704c8ff7703da0063027a02f200660201012f021904430398030b03;
// music[1448] = 256'h09036f04f105a20731075a06d70607073d074207ad06760740072905b9056106;
// music[1449] = 256'hd805ec06f0066407c4077b05a0050407fc045703570412059104ab033f035104;
// music[1450] = 256'hfc04be043305fd0440042504c50352034903ab032a040a0481036e038c038003;
// music[1451] = 256'h8d02d001de020403f702f502a301a202f40292029c039d022a0309027404f613;
// music[1452] = 256'h991c191aa41aca1a251aa51a9f1ac21a351bf21bbd1b201b1e1bd81a8a1aac1a;
// music[1453] = 256'h2c1a3f198f1952186a185719b317db191513bc0264008302bb007e0177003200;
// music[1454] = 256'hcd0089014403e5025b037a04bc03baffbbfcae001905b5077b093b09d709e809;
// music[1455] = 256'h1709a408e706210425022802d40157015301f60042001bfeb6fdeffebbfe0700;
// music[1456] = 256'h2001e600640254033b005cfd8afee301a9060507e7038804d4025c01f902f101;
// music[1457] = 256'h500369054c0699083509ff0a860c870d1d10090fc613101f12208b1ecf20621f;
// music[1458] = 256'h98214f2394206c2286202d237733b239fd369b377636a4359335c43435347233;
// music[1459] = 256'he532ab31f4306230472fc62d3e2c942b8b2abe29ec286f283a27a1258d274a1f;
// music[1460] = 256'hd20f500d790d940b580c750a410ac60bfe0bc10b4a0a430932087607ce07b907;
// music[1461] = 256'hc1069a07290b280c6e0be70bb60b890b540b550a27082e0882093b08e5086709;
// music[1462] = 256'hf906d7051206030765063b06d1064906a606340575050d052b0094008200ecff;
// music[1463] = 256'h9b010ff827efb6f0bdef5aee47eebdeb3bebf5ebc3eb13ec91eb4deb5bebeaea;
// music[1464] = 256'h2deb11eaeee95eea39e906ea7be953e925ea43e91bebfde8f4ec06fe6203e800;
// music[1465] = 256'h25034a02cf01cf029d02f002a603d4035503f7027103b905ac06980530051804;
// music[1466] = 256'h8903c1027d02fd011101fa0269fa07ec1cea61ea93e866e8dee86aeb56eb3fea;
// music[1467] = 256'hd9e9ade8a4e82be8dde7dbe705e7ade662e70be917ead9eac1ea14eabfe9b4e8;
// music[1468] = 256'h20e78ee584e603e8c8e76ee886e6eee464e63de656e648e752e77ee7b5e710e7;
// music[1469] = 256'h10e753e801e7b8e5e2e4f2e280e378e317e3cae3f0e3bae4e2e306e473e4cde2;
// music[1470] = 256'h1ae31ce3e6e221e30ee385e333e360e3dfe247e2c7e125e04de0f7df5fe073e0;
// music[1471] = 256'hfddf01e057db30e2edf390f7f4f57af7faf6fbf6ecf620f71ff778f65af625f6;
// music[1472] = 256'h02f6a8f513f6f8f56bf524f5cbf42df59ff406f514f5d9f55bf83cee40e021df;
// music[1473] = 256'h25dfc3dd99df77e028e0b9dfc2df7adfd1de08dfb7de26dedcdea0df55dfaae0;
// music[1474] = 256'h9ee273e2e1e33fe650e675e6bfe5bbe30be423e7bce89ee1a7d78ad95edfb4e0;
// music[1475] = 256'h0fe52fe8cbe80deb2bea1be9bfe8dbe664e5bde1cededadd61da4bd7b3d601d7;
// music[1476] = 256'hf7d632d73bd8ecd843daa0db8adc0cde44dfb7df7edf14e2b2e7e3e9dde814e9;
// music[1477] = 256'ha9e93ae99aea4cec3ced23f08bf106f49af775f70d0257149b1948190d1c481d;
// music[1478] = 256'h7b1eed1f5220e9204d21a8214322bc212a22d022f2213222a3221923b221e91f;
// music[1479] = 256'h0321851e401f881f5114ec12a218c31678187e196819af1ce41bfa1a2a1bd319;
// music[1480] = 256'h84191919651850181117ef157b17a718f417881753176c178f1754186e161e13;
// music[1481] = 256'h85136e10080c710c680be20ac40bd20b8d0c900c6e0cc90c820dce0dc40ddc0d;
// music[1482] = 256'he40b120b830b190a82081d069b04f604fd042105f4042004a90301043a04bc03;
// music[1483] = 256'h1203790262023f01f5ffa9ff08ffdbfe3dfecbfdddfd34fd16fe5cfe55fe3ffe;
// music[1484] = 256'he1fcea05fd147917c4158b175b16fa160f17b41426170512090661049705c204;
// music[1485] = 256'h2b04a80045ffdfff20006d00aaff6200130080003c015bf6acea28ec6fee52ed;
// music[1486] = 256'hdbed94ed95ed3aeefbed2cee49ee9bee1eef06ef9fef0cf00bf1b7f32cf430f4;
// music[1487] = 256'h87f6cef6bdf766fab8f9e4f999fa86f8e9f7daf7dbf765f8f2f705f84ff844f9;
// music[1488] = 256'h5bfad1fa3efcddfc0efe85fffcfdd6fc11fd00fd46fdd6fc71fb51fa63faaefb;
// music[1489] = 256'h85fcadfcd8fd49ffc6ff000089001e013c019801b6016f01e70117029102cd02;
// music[1490] = 256'ha90214030603fa03660350032b04f402910eb81e3c1f711e1420581f8520bc1f;
// music[1491] = 256'h4c1fd720a0209920f120f6206c21c9212d2145215721a52060203220ee20b220;
// music[1492] = 256'h0922ec2105162b0d7f0e990d270d100dd40b280c050c8e0b27090408de09cf09;
// music[1493] = 256'h8a09a909e109ef0b390ef10e7a0e740f7310a00fa3102f11a80d630b880cb50c;
// music[1494] = 256'h4d0cdd0c1f0d0d0d9e0cf20b390cd30c810c630cc40ce70c340de00be30afd0b;
// music[1495] = 256'h2b0b5d0ad60a6e0a940981075c079a08230860088308cf08b7096b09a1092b0a;
// music[1496] = 256'h4c0a360aca091b09b108e6083f080e081908e2077c086007e8077707cf05fc10;
// music[1497] = 256'h4e1d2d1d7a1c161da41c9f1c221cfa1b221b081b311b811a401a75196519bf19;
// music[1498] = 256'h2b195418bc177417c5162617c1169f17b017f10cc904ad05b8032c037603b401;
// music[1499] = 256'hf80112022702e5011d01340096ff6eff22fed4fe6000b9007e01e10025018b01;
// music[1500] = 256'hef007a00acfe1bfdaffc40fd0efd0ffc6cfc22fc2dfc7bfbc2fb80fc71fa7001;
// music[1501] = 256'h6b0c3f0d150c9c0c650d6f0ea50d600cb80baa0bf40a3c0a5e09e90704086108;
// music[1502] = 256'h7608a0086f083608fe075a08700818092d097208dc086c08a9074f07e506d105;
// music[1503] = 256'hb5047405b9044f056c042f045211bd1bd41a131b711a141a2b1ab119fd19c518;
// music[1504] = 256'h68181a18af17ab1759163416b516da162016c0153115b8146f15de13a016f115;
// music[1505] = 256'hee076e01db0281005effe2fe7bfe17fef5fdc9fd8dfc75fcb5fc06fd20fcbcfb;
// music[1506] = 256'ha5fdfbfd22feb9fddcfec8fe84f407eb66ea19e9e0e4c4e3d7e5d5e5d1e57fe6;
// music[1507] = 256'h2de67ae61fe642e5b6e4c4e45ee555e550e63fe6b5e4cfe420e5c3e423e459e3;
// music[1508] = 256'h4ee358e34ee3f3e3eae2eee0c1e1c0e119e161e194e04ee28ce337e36be476e3;
// music[1509] = 256'hbbe463e706e6b1e4ade3d1e312e48fe324e444e377e47ce41ce46ef0f0fa14f9;
// music[1510] = 256'h08f991f9b2f813fa9df9bbf817f916f959f9edf876f802f9f7f86cf88df796f6;
// music[1511] = 256'h41f75af725f79ff8d0f9a7fcbdf82bea43e5b3e720e578e5e9e597e4a4e5ece4;
// music[1512] = 256'h8be4aee4b7e380e430e4e2e204e5ace68de573e659e7f9e668e777e5f3e3fce4;
// music[1513] = 256'h9ce4bae311e4a3e52be693e571e506e55ae52ae5c0e46ee510e55ce530e6c1e5;
// music[1514] = 256'hefe499e4ede460e59ae5d1e421e497e2f9df4ce130e323e3e1e2d8e19ce202e4;
// music[1515] = 256'h59e4e3e447e5f5e519e67fe601e7f8e634e7bfe7d8e748e7cde731e7d7e64ce7;
// music[1516] = 256'h82e5c8e71ce768e78ff6f8fe99fc16fe13fef0fd99fee3fde9fd4efe57fe7afd;
// music[1517] = 256'hc6fd1efeccfdc8fd66fd9afc82fbf6fb47fb9afc1d00b3fecc0039fc7bec84e9;
// music[1518] = 256'h13ecabe99de977e97fe973e93de939e972e893e81de880e710e898e8a4e861e8;
// music[1519] = 256'he8e830e902ea46eba6e950e538e36ae5d2e659e747eac1ec67edc8ed5dee4ded;
// music[1520] = 256'h1fec1eec2eebe6eae6e9dee700e74be677e796e888e8e7e864e8bbe88ce86ee8;
// music[1521] = 256'h7bea70eb3bec91ebd9e92beec5f36df375f2ddf25cf171f19bf25ff21df427f6;
// music[1522] = 256'ha5f7f3f985fbb0fdfaff54018a0237049904d1053514a8292e32b43192312231;
// music[1523] = 256'haa30cb2f5f2fa12f5c2fe42e9f2d712c9b2ca62cf62b3d2bf029b92899288e28;
// music[1524] = 256'h31292328b1262829ea21f811fd0d0a0f4a0d150dd70b200c380b5609360abc08;
// music[1525] = 256'he5078b078e06bc0854086206b9070b09ed06e404bd056a0507068206cb04e705;
// music[1526] = 256'hda04cf030d0785070907c4075e07810779078d065a07cc0754051105ab05a205;
// music[1527] = 256'h130773065e065006a204b304a30351031804600487056a04cf0371032a03a305;
// music[1528] = 256'h2c0094f4e3f065f115f163f220f3e5f2adf237f2c0f2c4f1a1f104f238f1bdf3;
// music[1529] = 256'h47f284f5fb05020c380ab30bb30a310c750d2e0cf50ce40c570c550d780e720e;
// music[1530] = 256'h590f5e0f310f1b109f0fff1117138e12ac143c145f1633100101a3005b040803;
// music[1531] = 256'hb903c802ea010b011a004300efff78ff81ff4101f001750177017f011a01bbff;
// music[1532] = 256'hf000d60100014102af01e2004301e5008300940089027a033f03fa03bc035803;
// music[1533] = 256'h9b03520417031f027803bb03600444050306ed061606bd051205b6043c05d604;
// music[1534] = 256'h4d057b065206ac04760417053105bd06cc06ac079708b00792092e0a5e0adb0a;
// music[1535] = 256'h060a9a0bfc0a690ad70a8d0aad0cc60acc0ee31c8821fa1fba205c2031201420;
// music[1536] = 256'h0520bb2008218a20931e371cc71cf91d761d201eff1ea12004223420d520d320;
// music[1537] = 256'h5a20fc22c619fc0b810a450b440ca00d7b0cf90d350dfd0b850dda0bad0c590e;
// music[1538] = 256'hf90bcc0bbd0bb50aa30a5c095009b10a180ba00b3c0c1f0cb70b5a0b5c0b0c0b;
// music[1539] = 256'hbb0a8b0ba70bb20b0d0c180b180c600e040d23057afece029b077a09be0ebc10;
// music[1540] = 256'hdb1069111b108e0e030ccc0999079405e204d60283005dfe50fdecfda1feb6ff;
// music[1541] = 256'h4d019d021e03490493055306cc072e08ea08170cc81160136e11f41280100316;
// music[1542] = 256'h8f275f2c982c2e302f3179335d344c369338f639df3c2f3e174051412e421643;
// music[1543] = 256'h3243244554456745e7441d44e94397424543383a3b2e192fc72d892bee2c9b2b;
// music[1544] = 256'hdf29a92838277327df31ee3ca73b4d3a8d39a337d735c3329e327f32ae329b32;
// music[1545] = 256'h4f31fc316030402f642e742cf02b3029ae265d250c26cd280f2784235f20a91d;
// music[1546] = 256'hec1c8d1b561a101a9919ee186817e617eb1c011f0e1d1b1e2f1d6c1b481c571a;
// music[1547] = 256'hbb190719d91509152a1472139413cf12d511d610c50f440ee60de80cb80b480b;
// music[1548] = 256'h1f094a085207f6059d059b032b0a1817be19d91672174a17a315df14d8138613;
// music[1549] = 256'h9d137312df108a0fd60f7c0e6b0e4f101b0daa0c8a0411ee31e603e865e7f5e8;
// music[1550] = 256'hd0ddf8d0b5d193d173d0ccd1ead265d4c0d25cd1c9d23fd25ad1a0d108d179d0;
// music[1551] = 256'h2fcf65cdb0cd58cdedccd5ceb4ce2fcf7fd18bd023d0dad0a6d0e3d021d1c2d1;
// music[1552] = 256'h1ed093cee8cf1acf8ecdbeccf0cc9bcd3ecdbece3bd003d290d38bd139d1ffd0;
// music[1553] = 256'h62cf4fcfe6ce59cf1ad01cd062d0a2d0a4d0c8cfaecf8ad066d1a7d139d29bd3;
// music[1554] = 256'h2dd35ad319d456d47bd547d637d744d618d6a8d6cfd5a1d693d4bedcdfecdfed;
// music[1555] = 256'h6ded8fef98edffee8cee94eeafef50ef81f085f047f0d9f057f2adf373f348f3;
// music[1556] = 256'he8f287f3cff25bf3def3b5f315f41ae8bfddeedf16de77dd44deb2de29e106e1;
// music[1557] = 256'hfde226e3fce1e6e29ee198e153e055dec4dd6fddc8de10dffadf8de021e134e2;
// music[1558] = 256'h04e14ce1dfde6ddcb5de24de4cdfcbe1efdff3dd98dd0adeddde88dfbedf82e0;
// music[1559] = 256'h29e108e1fde16de137e105e286e181e140e122e255e17edeb5dfabdf19df7ee0;
// music[1560] = 256'h75dfbddf16e1f7e04de297e35ee3dce3ace476e44de413e4f6e444e625e6b4e6;
// music[1561] = 256'h28e7c9e763e6f2e46ef0dbfdc7fd11fc0efdd8fc83fdf9fc64fc2ffdf0fc8dfd;
// music[1562] = 256'h50fd0dfc7cfefaff81ff0200f7fe50ff36fff0fd44ff6dfe76002d01aff35fea;
// music[1563] = 256'hceebdfe986e981ea3eeaf1ed7af0baf046f007ef85ef22ee75ecc1ec4becc1ec;
// music[1564] = 256'hb3ecbbeccaed6beeb9ef61ef3df0e9f10ef040f0dbf08cef01f09df058f1ecef;
// music[1565] = 256'hbbec9fede3ed58ec0deea9eeebeeeaf08cf0c9f1c9f3d6f470f5daf230fdb711;
// music[1566] = 256'hf4153a131115a914c6146f15b1146b1488134013c514ec15b416f6172d181e18;
// music[1567] = 256'hd61766176718ac1951199e18a4180918301990183416e321672ef52c3f2dc12d;
// music[1568] = 256'hc92cc12e092ef02da72d972ce72c0c2db22ec22fa52fc02e842db82db02da32d;
// music[1569] = 256'h672e792f632ef62f342f791fae1552186e175c170618751ad51b9317ae18d019;
// music[1570] = 256'hff17ed17ea14b912ad135e14f81414158014ab14d214e1134a1470138a13b212;
// music[1571] = 256'h690fbe112410a3109e12a9fda9ede0ef8bed2cedd7ede8ed7eef51eee5efc4f0;
// music[1572] = 256'h8af02cf279f1e0f06bf1caf1d6f07eefa2ef66f01cf1fcf0b9f118f2fcf088f1;
// music[1573] = 256'h7cf116f15bf1e2f07cf148f2f1f111f2d8f15cf187f27ef200f2c6f37bf312f4;
// music[1574] = 256'hc9f3c7f2a9fe6d0a2f090b09780a5c099109c30b4a0d100ce10d6a1181103910;
// music[1575] = 256'h6c115a10c70e370fd90ffb0ea10ff60f8a0fdc100210eb0f7c10830f96123e13;
// music[1576] = 256'h2512fb140615a814d81224135f1505075df63bf4def43cf6e0f6f2f6ecf6e3f4;
// music[1577] = 256'hc3f546f544f480f690f66ef742f8dbf6aef776f70af504f5aaf5d3f424f57df4;
// music[1578] = 256'hd2f11af249f45ef437f337f3eef3ecf447f6b5f561f6baf7ddf6b3f610f555f4;
// music[1579] = 256'h3af64cf66cf668f5fdf308f3f1f2c0f5b8f5d3f5adf79af698f79ef71bf691f6;
// music[1580] = 256'hebf4dff424f755f66ff42af3fff2a1f56cf7c2f58ef56df7ecf799f640f87dfc;
// music[1581] = 256'h30fc41fdd8fce7f94b06e211c70ef410d817a61ac517f8103f0f51113e121713;
// music[1582] = 256'hc513021597147711cd124b16f9166019a217f9145315c8122617691354fffef8;
// music[1583] = 256'h74fa07f8c7f748f61af951fd1ef901f4f0f610fd51fd97fba3f902f431f129f5;
// music[1584] = 256'he5f891f91bf87ef2c7f2a9fa51f8fcf273f7d9fa13fa95fac0fc0301e70068f9;
// music[1585] = 256'h27f377f1c4f5d2f8a1f1c8ed35efe0f191f84bf779f1f8ef92ee22ef20f55f01;
// music[1586] = 256'hc3095407e5006801c508b107b9051a091308b104befd84fc94024d06b70ec816;
// music[1587] = 256'h631a0e189b12d314871d9c26ed1edf16e720a5200c292e40f746974903438733;
// music[1588] = 256'h733380386c3b0a3d203982376f39b63702368031142a4f2e72368a358831cc33;
// music[1589] = 256'h0739bc31a32a3428841b08137312b115d5164f13802056303a313a2c80222b21;
// music[1590] = 256'h3129d732af3a1238923099284727ad2ee430e832b036ae3681355930092c1d2b;
// music[1591] = 256'h2d28d82a2c32cc36e839ee32b228602e3b30361c430a090ecc1a9223c0298728;
// music[1592] = 256'ha023f3227d217a207619410e1c0e590ebd053cfd56fefd040f06c0085e0772fa;
// music[1593] = 256'h70f544f890f914ffd70585079409dd0ed40c1b056e06650d6113411b261e981e;
// music[1594] = 256'hfa2a9636143a5f3edf3c293d693fbd380f3b98432e46914825466c458e4d2851;
// music[1595] = 256'hc246a8371136f43e2d441f4622480747ed3f7432f123e21e29216025d0293628;
// music[1596] = 256'h8e28472b73240b1ebe22902b52306b307027fb1fe729ec2ddd265726c127a62c;
// music[1597] = 256'h662dfd29f727ca1b42189720cd1bc015a0185c1ec0296531012af8209b1a7b12;
// music[1598] = 256'ha8120a17a31b9522a8202b1a21180d18ab16f114b01974218821db1b29181317;
// music[1599] = 256'he6190e1ba61352146919af18481c721a96163b18af187a1a69141c0e840b5503;
// music[1600] = 256'h650964170a189114111b1e2ae62f9f2acb26a8276c2bd42e772f4425ce174b17;
// music[1601] = 256'h891ccd208f285c2e162cc42bf62b6820911aaf222527062a262f42252611ce06;
// music[1602] = 256'h34002501030e5c105808bc0137034c0ab40a670c590c3506f5073d0892020f00;
// music[1603] = 256'h650047039404e801720127052f06c20199fb88f8acfbb0f977f59401090cbc04;
// music[1604] = 256'h2300eb013004f30592fca2f5e1fcb5010503d402560060fd73fb3efdc3f48ceb;
// music[1605] = 256'h57f0eef370fb8606f108ff010ef623f6d7fd3100affe98fd67ffb4f946f400f7;
// music[1606] = 256'h7df80affe303d8ff13fb55f7c1f354ee6af3a50b6d1e731cc915dc11d50b800d;
// music[1607] = 256'ha6147416d315f014d11524150411de0e5a0c240bf00f3b17b615eb0dba0c9511;
// music[1608] = 256'h421a521b1d0d65fd5df246ee58f3befc22fa71ef12f849010efc16ff9f0350fc;
// music[1609] = 256'hc6f0e4f3dffc5af142ec9af890fbcefcf3fd9efaf5fd87fd8af71ff8e9f9a6fb;
// music[1610] = 256'haef734ec31eee2f529f7b9fc5ffc05f712f65cef53edd7f80a0214015efc11f9;
// music[1611] = 256'hd6f6d2fbb103e8fffbfdf209e0143619681d041a8206fdf9bd0563136a17df14;
// music[1612] = 256'h5a0bb5091911960e540772085d077905f30d5d0f240479fe6a06b916181f1e23;
// music[1613] = 256'h6229ae231e1c941cd719b3160e1b3e223c200418f8151715e7133d1c8225a923;
// music[1614] = 256'he11f351bf313d411d10f9a0541f309eedef82ef3fced59f87afb9200a507a904;
// music[1615] = 256'had004000fdfe62f7ccf2f9f250f083f443fd9cfc4bf6f2ed2fe3c7e533eeb7e5;
// music[1616] = 256'h8be0a7e361e23ce5b0e5cbe121dce1d596d55ed7f8d88ccc6fbae9ba82bc11bd;
// music[1617] = 256'h6cbedbb550b4b6ba3fbb14b5b7af48b26ab427b823bec2ba6fb4beb1e6b126b6;
// music[1618] = 256'h62b976b363a75dab85beffc33cbdb9b9e2b8c3b6a2b272b425b85eb978bf71bf;
// music[1619] = 256'h33bfc2cb75ce66c847ce1ad7bed962dd39df42d549cfbfd7b4d999d5a3d87ddd;
// music[1620] = 256'hf2dc4ed79ed88cdca7d70ddc10e6e2e487e0acd4f5c73bc79ac601c774ca99cd;
// music[1621] = 256'h65cf3fcd77d166d623d38dd233d1cecb1ccd77d57ed3d8cd06d6c3d706d2bfd1;
// music[1622] = 256'h67cf9fd6a8e225e033d52fd0afd608dbe8d589d1b3d28cd57fd737db1cdb35d6;
// music[1623] = 256'haad4b6d456d1a2d077d964da60d8a3df35d698cc94d227d074d566e2b5e167df;
// music[1624] = 256'h2ae01cd953d2e2d993dffcddeee423e623de07ddeee168e5c1e360e245e3bfe5;
// music[1625] = 256'h7ce8c1e141dfa1ee12fb17fcb1fe90068e0b3105a3fc3afc0800d7047a06bb06;
// music[1626] = 256'h5506ba012d0185fffbfe3708a1073f0154019b01ca034efdbef30df28aecb3eb;
// music[1627] = 256'ha8ec3ae478e6b6f4c3faedf51ef0c5ed6eed9bf1cdf487f081ebeaeacbeec3ef;
// music[1628] = 256'h55ecf3ede4ee65e8b9e06edf7be5d5eac9efe6f1f3ee0df0f2ef42ec25eb33ee;
// music[1629] = 256'hf9f3fef010ebc8e9bce6e5e5b3e47ae449ebdcf142f52df4e3ebfbe1cadfccde;
// music[1630] = 256'h8ddbdae230ec41f03ef1acebede567e3a9e758e923e076e1f8eb4cf032ee57ed;
// music[1631] = 256'h90efe0e9bfe604eb78ed75f628022b0b8f0eac0c710d850bb40a80089cfd37fe;
// music[1632] = 256'h5407dc0a021217167e115e0c1c01a6f921023a0a310b450ca70e560854fc7dff;
// music[1633] = 256'hb106db08520aba049806aa0bc4052806500f21129e095c037a07830a50056700;
// music[1634] = 256'hd007690c120afa0cb409cb0506045dfff904d40a4f0c170f290d0f0bee06f5fa;
// music[1635] = 256'h35f42cfab200e1052309b0ff35fbc902880277007803dffe43f60df8f9fe1c02;
// music[1636] = 256'h0a05e10263f822f145f697fd3400f0034701eafa35fc74fe32ff0efe08fb9ef6;
// music[1637] = 256'hd5f6840101023af7e3f7d9f652f3980b9b23c119dc156d19b1115d1757185d0f;
// music[1638] = 256'he7133f178618e618b012f20ad000e6fe700294fd61f952fdb2fea3fe8304d8f7;
// music[1639] = 256'h62def9de7be8cae727e612e4ede5cfe759e29dde7be55bf066f597f912fc2ff8;
// music[1640] = 256'h9ff10de880e43ee9d9e70ce9e5f247f5cff2d3f393f25ceb63e344e523eb37eb;
// music[1641] = 256'h4fed9df0f6eaede4f4e932eae7e000e389e9d4e8cbe587e4cce968ee1bf180ef;
// music[1642] = 256'h3ae52de4f5e78ce524e307e1a3e212e5c4ec91f272e406dff8e629e683ec54f4;
// music[1643] = 256'hdef0dded07ed8fecf7e726e508e999e7a5f029067a073f002907020e2e0c1a05;
// music[1644] = 256'hc5fc68fb78ffe801340644091a07ec086f0a2009c60c8c0be6ffecf5dcfba307;
// music[1645] = 256'he1fe6cf004ec8ee275e353f217f3fdf1d0f492eabbe737efdbed9beda4f2cdf8;
// music[1646] = 256'he7f747ebc5e7ceec9cee1bf462f7aef395ee39eb7cecafee48ef3aec1be634ea;
// music[1647] = 256'h72f52bf374ea21ed96ede9e2b6dfdfe632ee82f292eeece82ce95be781e310e6;
// music[1648] = 256'hc3ee96ee8fe7cbea45eabce66eedfaeb6fe4b1e05be373e9d8e18de183efb2ef;
// music[1649] = 256'h34ecafea32e853ed8ef07fee75edaeea54eb3cf9020b1e114a0fa910f2109f05;
// music[1650] = 256'h7ffce3fe7d0022006f01170bc311050959068507d30985124a11280edc066500;
// music[1651] = 256'hec0723fd5eeb16ea0ce8eeefe6f768f192f05dee9aeb49f0a7e826e65af33bf5;
// music[1652] = 256'hd3f690fe5afc48f64df07deba1e997ef42f8e8f2f7ed71f5b9fdceff8cf9f3f4;
// music[1653] = 256'h0ff742fad4f526ee33f0b3f2d0f496f189e6e9eadfee81eac0eee9f41ef911ec;
// music[1654] = 256'h02e015eed3f283f0d5f322ef21f7e7ff1cf86802c514390fde09fe0cf7095f0b;
// music[1655] = 256'h661254181a184714501a7b1cbe1b4a21e3233137b64b35438d3bbf425749cd45;
// music[1656] = 256'h2e410048914b6e49a448a441b030f6255632c73fa140e8428b45e4436e3ab739;
// music[1657] = 256'ha844f3363d1d90186215a10d5810ac0eec078009e1067108f90d7c069607910f;
// music[1658] = 256'h160d480a2109100dcc13e7142716a01743127d0e32135b1227129219b41c1723;
// music[1659] = 256'h43273e23ca1f43184516ed1e5328842ba22a1c2c1029352a0e2c9c224227092c;
// music[1660] = 256'hf11eab1b671e1c1a32179c170719c41a561b0d1cb4221b23461aac1ca121db1c;
// music[1661] = 256'hbc190d1baf1d2a24912b1e2c562d402b1420a12a6f3fc441be455147a640893c;
// music[1662] = 256'h5b38d33d8942f13cb03cb040ff45fb45053f873e2a3d23356f35723aa337053b;
// music[1663] = 256'h053d4a262b13f515c81de7203519d4168b24f227921ad017bc1f2c20b7222323;
// music[1664] = 256'h611f412490225e1d441b1817f81b0f1bbd14bf174916f215921b2d1cc919ad18;
// music[1665] = 256'h2717be15851c481c800e430fce126c0970055b05ed090414fd14a80f4b0c220c;
// music[1666] = 256'h8a0d260b3b0202006d0c800b47014108320bdf02eafee1fe83ffaa0240099504;
// music[1667] = 256'h3c017d046afe2705b10aa1044809ec07cf104f22fe1dcb1bdf1f8a1e041efa1f;
// music[1668] = 256'h101f171cb820b91d1617951c1b1b32163919621b0719191bda1bb012aa16cb15;
// music[1669] = 256'hb2001802290a8606da0963029ef412f334f568fb190097022f09930a230ae305;
// music[1670] = 256'hdafdad0397072307a009e4034d08c60e0e07770469017800240c0112730a2308;
// music[1671] = 256'h7c0a3e07660a2e0846fedcfef7fd3f04e5093e033807cb0340fafdffdefdb2f6;
// music[1672] = 256'h39f9a4fec2036d0199fb4efc5ffbecfcc8fe12fa65015e070003c4002af6dbf6;
// music[1673] = 256'hbcfc90f62ffe85023afe9f027205e60e251e401f43153e18541fd717c31a2a21;
// music[1674] = 256'h4e1d231f951b0416a7199d1ae919471b901a8115e5103a14021e0a1ee50bc3fb;
// music[1675] = 256'h32faf8f91bf70bfacd020809900619028904b8053104dd08600d0e090708d311;
// music[1676] = 256'hc8138a0de60a470d501a5d206221d725331ca61ae320971bcd1a901b98207721;
// music[1677] = 256'h331aff1da91acb121111740d7d1480141b0cb512cb161713a60d890620074507;
// music[1678] = 256'h620ab913610fee091c103b0fc505a900ae05e20a5b09670ac50f730d1e048205;
// music[1679] = 256'h5304f8f7fff775f91500fd10a311310fa411ca13251a8219941521179f1dfb1c;
// music[1680] = 256'h1a18291ce5182313d5112e0e8b08a9feb804f30be8038a0469fc5eec9ee504df;
// music[1681] = 256'heade54e217e101df73dc5bd9aad954d9e0d257d5e3d38cc90ec717bce1b54dba;
// music[1682] = 256'hfab71dc06cc47fbd2abeb1be48bc58bc46c016c323c43cc4f0bd0abc52bdbbbc;
// music[1683] = 256'h84bf27bda4b81fbb4ac064bff8b925b56bb089b4e8b88bb8fdbd6abae4b6bfb9;
// music[1684] = 256'h5bb5aeba2dc1b1bbeab617b534bbe8bdbfbc4ec347c0a1bde9c6b1c4c2bd7ec0;
// music[1685] = 256'hc3be62c128d47ddf9ee17ce301e2b7e7f0e67bdf35e694eab0e59ae09ddd03df;
// music[1686] = 256'h71e04ee3c3e725ebc8e8ede8b6ecd5ea09f249ede0d6a6d2e2cd71c99acd0acd;
// music[1687] = 256'h69d129d0cdcf0cd69dd596d6efd4cfd431d566d499da1bd9cad815dbc3d895dc;
// music[1688] = 256'h5ddc1cdc7cdeeada18dc18e126e388df50e04ce88fe5f7dfb5e022de9cdf32e4;
// music[1689] = 256'h4be17be1e0e473e32be66ce48add0ee17be589e3bee1b3e084dc9dd89eda91dd;
// music[1690] = 256'h8be0fade9bde09e3a3e1f8e054dcb3dba7e592dff5db96e1c5e0c4e4dfe456e8;
// music[1691] = 256'hbff852007afb84fcce068506cc016d0081fd3603cc04db01f7032c030b0221fe;
// music[1692] = 256'h9efcbbfe5f00ad04dd0120019cfa52e67fe1dee276defbe2e4e680e2d0e162e7;
// music[1693] = 256'h6ae573e3eae790e597e62decb1e6cfe5e3efbfed01e248e0eae5daee28f69cf5;
// music[1694] = 256'hc9f28feecaea40ed9bf1e9efadeb33ed75eebdedadecf1e7e0e6cdeb50ebd0e1;
// music[1695] = 256'hfbe0d8e9b8eb50f1ccf314ea3fea21e9c0dedadf29e60ce506e116e310e909e5;
// music[1696] = 256'h02df33e565e9c8e8a1eb2de8bce5cee9c4e8b9e64fe404e6cbf43e00ab008603;
// music[1697] = 256'hc4097b09250461022505530552024d05a20ab009c8060808e70a70083d0f8221;
// music[1698] = 256'h12274925531f270e1d0188faddf883002608c909320b3c0703fcd1fcc9003efb;
// music[1699] = 256'h11fe7101e9028a09db079a0462017bfca7fd18fb77fd5d0741061005e1093b0a;
// music[1700] = 256'h37083c0565028c038e06770624038200a100150426079d07430a480b16031dfb;
// music[1701] = 256'h68fecf02fbfe94fd880058fd65fb9bffa7fd7bfca50287014efea2fe52fd79fe;
// music[1702] = 256'h25fb66f99cff5cfd1dfdaf006afabefa6c05260e67115712fa15c61433108412;
// music[1703] = 256'hf9173a1726127216231a2a0d21fe74f828f978fb7900cf0722067900faf8f9ea;
// music[1704] = 256'hd8e4d2e504e7efe8ffe519e4cbe5a0e64ae602e778e997e2c1de0eea39ebb5e4;
// music[1705] = 256'hd5e793e664ddb6ddb0e773e92ee60fe844ea08ed9becfae8c7ec62edc7e55ee6;
// music[1706] = 256'h0ce938e758eba7ea50e6e8eb22f0daef4aed1ce854e738eb1cede3e85eec9cf0;
// music[1707] = 256'hf8e7cbe558e631e8cbeb9ae4e4e361e61ee88cecf9e8e2ea15e6d2dc8be21ee4;
// music[1708] = 256'h85e8f9eb85e47fec9cfb6c00750359089b0414fe41016c038e060709e403a203;
// music[1709] = 256'h7d03fa03100a7f0bd60348fc4e00f801ad03230714f623ecabef0ce781e415e8;
// music[1710] = 256'h1be552e09ae51ff24ceea5e978ebc0e8e9f0c6f182e80debfbec74ed56edcdec;
// music[1711] = 256'h30ed84e822ee58f430ef3bf0bbef42ee5cf3c1f0e8ea02ee77f0c6ed1df0e9f0;
// music[1712] = 256'h4ceb3aec03f055f139f396f4f5f3adf010ef6df07ff12bf0baed51ee0ff2bff3;
// music[1713] = 256'ha3ecc8ebb3f3a2eeaeeb3def92eb34ea6de8cce7aaea84ebc8eb28e8d1f15507;
// music[1714] = 256'hbd095f007b010d0af90b280917074e012704890bad07e806da074a04f60a760d;
// music[1715] = 256'ha505f708460d25090701f8f1f8ebd8f02af201f21ef0fcedd3ed9ced18f000f3;
// music[1716] = 256'hb1f1f3eeb8f083efd8ead7eedfeed2e652ea44f4cbf4adef94ec66ed39f41af6;
// music[1717] = 256'h7bf23cfb4eff8ef493f04eeeb2ea8fee9ff3f6f6d0f822fcd4ff9afd20fa26f9;
// music[1718] = 256'h0ffa98f996f594f395f28ff057eedfec97eecaecc2e9fded48f630feacfe5bfc;
// music[1719] = 256'h04fd83f545ec74ef9dfa3a0168fd14f8e904f1246032d0287e2c1133c02fe52f;
// music[1720] = 256'hef333b39fe39cb3c36454644753eb53db53fa53d003bba418842e33fb3496e41;
// music[1721] = 256'ha927e423e527212984296818761348202d225329b32be825c729ad248b215527;
// music[1722] = 256'h52216f176111ce119013130f630dbc105c12ad10e00c3e058003330ba609d607;
// music[1723] = 256'h0e11f4153e127f0cad0d8d14bc19131beb1bb9216c212321832792257e28742b;
// music[1724] = 256'hb526fc29eb2720290c2fc5298630c233eb2bbd327a33c830b8376739ff372a2e;
// music[1725] = 256'hb31f241dcd23e6323740e03f173f9f4370423b3f2c40ad3fa13e5c3c6e3ae13f;
// music[1726] = 256'h384253417c45a542ca3eb145be45f24325468233d821f925b2238822e0275b23;
// music[1727] = 256'h832290261824e62210283029c722671f341f531e441eb323ad26051e30205926;
// music[1728] = 256'ha2219925b723931c8b2178228d24422606229722f01d4718391c39203f1d6e17;
// music[1729] = 256'h211ae71ddb19a516791aed21b51f6719ab19ab1c7122181f2d19c91ea21c2815;
// music[1730] = 256'h45138513c717cb16af1197113612f514fb199f17830c720a69183e240d246920;
// music[1731] = 256'h0520c02148245024d824ef2795231e1f37206022b5288429e4249a20e21a7b1b;
// music[1732] = 256'hb3205b23cc19ed066f01e407960a8606bc04f80473fef9f9c8fe130461014402;
// music[1733] = 256'h400872027003480722fdf9fe650473feedfe980355045d021303920529026cfe;
// music[1734] = 256'hab04de0942063006c002b0fbd501b205c1004601c00456044d029500b0000606;
// music[1735] = 256'hea04bafd2b02b60ab60e500957009c064f0c95041902e1047102e804f2090d05;
// music[1736] = 256'h0c036f05b2085d0a7f027a08ae151d1863209820b717db150317fc1b521bb91b;
// music[1737] = 256'h7d214d1e791c161ce51b54225b1fdc19ef1aab194920331e9504bbf71bf9bdfa;
// music[1738] = 256'h660271ff83fb9b023503330419046fffc600540067fe200034046004dffcd000;
// music[1739] = 256'h5406d1fb8bfc6c06080296fda0ff26ff5f005d037305da067303bf0033022703;
// music[1740] = 256'h5c05cb02bbfd5d004b023dffdffde1ff6cff45ff3907e70a990c9911030b2908;
// music[1741] = 256'hf6109e0f090dfd163f1e421cba190619001d411ef719eb1e951f201d5d29d22c;
// music[1742] = 256'h012a142ff729a122e5241b28ad2a872cdc2ac4293d2bfc28ca28fd2f9131192c;
// music[1743] = 256'h6a28a628712bf2249d115f074c08b2063009900b6a075905b20277ff92fd10f9;
// music[1744] = 256'h11f31ef1d1f510fa9bf9bef825fb2efc5ef628f525fc3301560021feedfb23f7;
// music[1745] = 256'h38f74df7d3f457f653f230f5dcfa7ff187eb4decffefc2ee07e67ee8a5e9aee4;
// music[1746] = 256'hdbe394e2dfe1f3de56ddf6dd42e002e353dda1d742ce2ac21fc225c114becabc;
// music[1747] = 256'hdeba15bd3dbf5cc133bc36b5e4c4b9d621d8a6dab4db30d628d038cb3ad197d9;
// music[1748] = 256'hfdd4c6d2a5d6f0d3dbd036d1d2d23bda50dd07d6b6d764d97bc9e6bdf9be7cbd;
// music[1749] = 256'h80b98abcfcc075be26c170c30abe47c015c4a5c486c6b8c24cc021c489c422c3;
// music[1750] = 256'h7bc538c50dc50dc8a6c6b4c7a2c9a3c4c0c45fc9c5c92fc7f4c7c0cb0ec9f1c8;
// music[1751] = 256'h4bce36ce6cd4e3da9ad187ca44cc43ceddd02ed04dcf36cfd1cf90d6e1dacadd;
// music[1752] = 256'h3de4dbe458dea5d509d6dfdb1cd9c4d82fdc85d9dadc26e296da4fdd5cef0af6;
// music[1753] = 256'h16f907f9d8f365f60df5c3f67efafcf3f3f026f07ef77ffc2cf6f0fc92fc08f6;
// music[1754] = 256'h40fc51fc7cff15fcf4e5f5dd8adfe6db48dee0e1c9e132e248e018e214e4bcdd;
// music[1755] = 256'h4cdffde495e2eae3a4e257dbbcdc1ee327e2e8e4a8ed74e73fe48ceb61e437e4;
// music[1756] = 256'h38ec48e5dbdf9ae0b9e229e629e65de656e743e860e80de814e9f8e800e86de3;
// music[1757] = 256'hf3e0c9e5c9e62fe517e62fe79aea38eed0ebdee62bec16f3c6f17ff4d5f667f6;
// music[1758] = 256'hd3f2d2e967e991e62fea3e045b0e15099e08e4079e0cf50acc04cb057b02d801;
// music[1759] = 256'h68074d085c048b0397067b048d028e018f00730493fa36ebf6ebe6eb05ea1beb;
// music[1760] = 256'h5ae71de74feb89eec9eacde39ce90cef22ee68ef3ceb8eeafbe99ae72fef5aec;
// music[1761] = 256'h39e7acefcaf073edb1eb8de952ebfeebc0ec3aeed3ea0ae7cceaa2ef30efeeec;
// music[1762] = 256'hbfe849eab4ef8eee76ef2aed89e73af00ff53ceab2ead1f2d3f134f51e000008;
// music[1763] = 256'hb609240af60bce0a270dbb096304400d510add006f01e106551bb0222e1db323;
// music[1764] = 256'he921c11da31d4419c01a261e5e1d411bc41cb01caa17a21588188d1db01cbd19;
// music[1765] = 256'h9816da0a8701fefc06fe0c041a0030fb49fb7bf93bfd3b014fff73ffa2ff6702;
// music[1766] = 256'h6104edfaf2fb4f02a9fb45fe6c01db016503a8f844fdcd03adfa8100a30042f9;
// music[1767] = 256'h1cfdbaf8fcf460faa1fa7ffb10ff2dfc41fa06fdc6fb7ffd0101150052ff30fb;
// music[1768] = 256'h94f682f4d1f6e3fcc3f43ee9f6e93ae7ace374e75beb30ed8bed0dee02efa2ee;
// music[1769] = 256'h15e70be5ccfc960c420312039b063907bb0a5803e3fe1d030b02af0262047705;
// music[1770] = 256'h9c09a6075103fc0345fe1cfefe0722fbd8e4b5e1dce5afebb2ed09ec44ea81e5;
// music[1771] = 256'h7fe45fe6e0eaaaeb33e4c4e403ebd2ed95e95de4c5e5c8e3b3e52deb77ea9fea;
// music[1772] = 256'h5de9e4e9c5e941e8a3ec91ede0ecdee700e3a4e7d6e45ae5caed39ea17e85bed;
// music[1773] = 256'h69ee94ecf6eb60e91ae750ebd2ed76ebb1e9faeb1ff2a9f0ceebcaeddaf147f1;
// music[1774] = 256'h3dec4aec63eca1e858ecc9f164f1c8f0c4f87a035e07350dbf10800ef30a4f05;
// music[1775] = 256'h1a0594032105910eed0bd009210d780cdb0d1a06b6008708d60ba408fcf81fe7;
// music[1776] = 256'hcee93af266eee9e7aceab1eb59e766e62ee68dea24ed75ed4cf305edf5e6f7ea;
// music[1777] = 256'h1ce774e83eefd4ef5fed42e95eec40f084ed22eb6cecd5f032ed13eaf8f011f1;
// music[1778] = 256'hc7ed31ed0feaace961eae1e878e86dea3fec93eca9ecadea2ceab2f0a5f2c8ec;
// music[1779] = 256'hafee05f150ecf5efeef365f1a9f3daf487f265f3e4f416f563f39fef15f6c408;
// music[1780] = 256'h720e950965082a052308990bdd09990c870a430adf0d5407d004030d580cce05;
// music[1781] = 256'h750dd3116b0dde116706eeef07ec2beee6ee5eeca9ed51f585f195eba1ed2cf1;
// music[1782] = 256'h84f212ecc5e751eb98ed2cf141f78cf7f1f4f6f227f155f51af74aef90ebbaed;
// music[1783] = 256'h30f0b6f093ecc2ec44f2b6efa6eb9aefd8f36ff5b9f1f4ee4af4eef2c6f2eff7;
// music[1784] = 256'heaef61ec60fadc056e04c8017a0422055f0e41189817f11e1e20751cf6228121;
// music[1785] = 256'hcd207324ee28b52de626ab34f14d1a49d643ac45ec421d49ee4a02443b45734a;
// music[1786] = 256'h36492949be4347326e31de3c76426248b447d348e845962fd2201821f521551f;
// music[1787] = 256'h921ddc1bd411080b200a8f0a610ee80bf409c40a65097f0b670c420efe120114;
// music[1788] = 256'h14157617e013500e4313e618af154c18b922c322541d9422532359234a2ab726;
// music[1789] = 256'h80285a2c6e29a42ff12ded2b71300330fd332833fd345b3c933c9042093d8b26;
// music[1790] = 256'h5e1c49226828ea24a222c82597262226e3244029b430cd34dd3b1f441c487d48;
// music[1791] = 256'h5b456f41ee3fb33f0342ea452b4481412042c941eb412f41cb40673f733a3d3f;
// music[1792] = 256'h4e43c9314a2046216428ab28da20d71fb527f6276820bb1d512184205c200d25;
// music[1793] = 256'h78224b218321ac1cd91ca11c8b1f2423dd1bab1a8b1cc3181c188c16f118ff21;
// music[1794] = 256'h422007178f185619bd14e018b61a051a871b4f168313b311aa0e250fad0fd013;
// music[1795] = 256'h34145812d616971684157917ee157d15a114210fcf0dec10d40e140d3e0f6b0c;
// music[1796] = 256'hf2070710a8227229e326fe25b225b92aa025f01f6527842442264f27321cc520;
// music[1797] = 256'h9623cd2101240122ff255e22a01dce1c4010550acb0412ff1603fc0068fc6bfa;
// music[1798] = 256'h07ffcd040201a0ff2d00a203f0044dffc502ff07ef0435005c0382082d026700;
// music[1799] = 256'h8c04ac03340378033d04e700e6016a04bcfe960095015ffde8fcd9fc78022002;
// music[1800] = 256'hb0febefe7cfa4bfe93022d02d40599050606b107da08930b050b45080b03d9ff;
// music[1801] = 256'hdb05780a34040700f700df0162080e06b4094e1f711f551c17205d199b1f761e;
// music[1802] = 256'h1b18e922cf1e7316b918151bd21c1317b619b321641be918a41ece1b9b0c2600;
// music[1803] = 256'h3e0066ff5dff2904580145ff0602e9fda6fb04007bffdffcbdfde0fb23fa10fe;
// music[1804] = 256'haafe9bfe9705c4059cff6cffbb003c05cc08ed025100cd000ffd4ffe90ff24fc;
// music[1805] = 256'h11fdedfe8502b008f107ef06b50544feb3fa66fbe6006d059f00d103a1098408;
// music[1806] = 256'hbd0a1a08870e9c1f2f1dcf181a20c520171e061f4d1d8115ec13d317d6171622;
// music[1807] = 256'h402e032c4b2aca2e5432512fc929d62bef2d5328d220bf2023264f271328e227;
// music[1808] = 256'h2f24392306234623551cf70aab03380626055402c901c90224fe7bf5fcf1bdf6;
// music[1809] = 256'h09fbe7f73bfa87f939f129f6bcfbf1fd44020a008effe9fb1df9ebfd8bfa43f7;
// music[1810] = 256'hc1f625f466f4acf379f1dfefccef1deb24e627ead9e7e3e2d5e245df90ddddde;
// music[1811] = 256'h45dc57d995ddf7dc98d750dddeda7ed670da6ecc40c2c1c84ec527c1a7c1afbd;
// music[1812] = 256'h2dbc5abca9bb11bb1dba00c672d5efd31fd10fd4d6d55dd472d3fad8e4d5ffd2;
// music[1813] = 256'h68d8ebd5fbd848dd9cdab8dcefde64dd98d820db70d86ec17aba00c5e2c641c5;
// music[1814] = 256'h4dc41ec018be22c267c16bc1efc4bec1afc40ac740c5f0c66ac2fdbda4bb88be;
// music[1815] = 256'h4ec7aac73bc854cb8dcdd0cddbc9eecac0cdddd006d1b7ca9fcbd7cfc0d1b6d2;
// music[1816] = 256'h58cedbcb02d2b1d7dad2e1cffdd025cdf2d0fdd507d2edd05cd212d6bfd92bd6;
// music[1817] = 256'h34d495d96edc15db8adb85d982d605d9cfdb6adc18db35deb7eb4cf51cf594f6;
// music[1818] = 256'hb6fb3afe0cfb87f804fbe2fb4ef7e8f536fbc8f77bf2a1fa13fb46f737fcc2f9;
// music[1819] = 256'h4af927f645e4a1df0ae63ee409e11ce254e3b4dfe1dd96dfc5e0bae207e290e1;
// music[1820] = 256'h62e06edee8e1d8e486e421e27de043e3a1e3c8e1e4e49beacfe764e059dfede1;
// music[1821] = 256'hf1e76ae955e7a1e91ee4b4e2cfe743e5e3e80aea8de640ea9ee9fdea91eb69e5;
// music[1822] = 256'hade656e66ae589e94ce6a6e5a0ec30f02af062ec50e9b7e995eac5ec0bedefed;
// music[1823] = 256'hb2ece2e8d8f6e1054301fa008b043803b605a4056c047b09230c1f06e3045108;
// music[1824] = 256'h5903ea032b070405e9073805b304ea03bef0c2e877ec68e9f3ea50eba4e9d1e8;
// music[1825] = 256'h51e5a3e7ffe945e7eee5bce35ee1dae39ce8d4eaede94de9b8e97be80de91cee;
// music[1826] = 256'h00f065ecfee9dde9c0e6f8e355e7d6eb24eb4ee860ebb6ec84e714e8fae7a2e7;
// music[1827] = 256'hd3ec33ed53ee4eec5ee821ed4cec68ec71eed9e845e9a7e81eeb82fba6059904;
// music[1828] = 256'h360248017601c3037805e603e804e5015c041e14f5173f192f212b1f481d8f1e;
// music[1829] = 256'hec1e791f591f1023cb207f1a6f1bf31b421ab619281b421b7f1a551bd8100a02;
// music[1830] = 256'ha9fd66fe300155ff45fba9fb0ef85af653fd4700f9fdf9fe29fc2ef924fde9f9;
// music[1831] = 256'hcef8e7fd80fcfbffbbff18f9acfaf8f9bafab3fefafda2fc55fadbf935fadafb;
// music[1832] = 256'h1e000b0045ff95fb72f8f8fdadffeafd4cffb6fbe1f8dafc37fd9cfbaafd2dfe;
// music[1833] = 256'he4fe58fd49fa7ef807eda3e5ffeddfeed5e6bae8a5ed0ce854e4f8e52ae660f2;
// music[1834] = 256'hea00e7020202e3fecb00c4077406c703cc03ea031f0552062e04d7fd2cff4406;
// music[1835] = 256'h3807d3064307a40773fe53ea97e532edabedf8ec6feb32e7ace785ea52e96eea;
// music[1836] = 256'h20ed8fe90beb70ed0de836e690e559e7cee887e55deab7ec18e898e6a4e6c8ea;
// music[1837] = 256'ha0ebdbe8f3e97aeb69eab2e608e832e891e321e5b8e67beaf6eccbe77ae779e6;
// music[1838] = 256'h07e282e3c4e7b4e8a4e559e7c9ea4ceaaeec1bf04af0feeeabedbded0bf1cff2;
// music[1839] = 256'h20eddce9feef76f42af063f51607aa09ec04d9079508970a490c1b0ceb0dfe0e;
// music[1840] = 256'hc30e930ba90dc40eef06c204c90511078108070a190c32fc7fedfdf04af08bf1;
// music[1841] = 256'h96f32feebced2def6eeea4ec88ecfeec6cea48eadee96beb02ed14e93aecb3ee;
// music[1842] = 256'h2debc1ec28ec20ec31ed19e8a6e84eeef6ed3decc7eccbed98ef1deee5e907ed;
// music[1843] = 256'h3bf2deef98ed5aed9aeb42ed9aef9ded1bec53edaaeee2ed8aebdeecfaf0b0ef;
// music[1844] = 256'hc5eb32eeefed2ae983ebfcedbbef19f24ff0e8f23ff01defb5009a0c330d150c;
// music[1845] = 256'hf208d70ae40c750dec0d710e8b0e210c980ff610a40e510f600ae70a980cda06;
// music[1846] = 256'h9f0aaf07d4f6aff01ef169f054f4d1f366efccf133f29eefbdf0f0ef04f1edef;
// music[1847] = 256'h91e7f3e7afee6ef15ff6cdf7d4f32cf7cafcdaf95df624f9c4f7e7f025f09ef0;
// music[1848] = 256'h1ef0cbf049ee26ee4eeed0ef0ff4def140f38df35cf04bf59df4a9f003f0a9f1;
// music[1849] = 256'h4dfc0d0162fef2fd45fe5afd5bfa93038413f71731180a172219ea1f38211725;
// music[1850] = 256'h2f2aaa272833f147ca499947f3473744b048234af7447b44274445481b507c4e;
// music[1851] = 256'h303f6f34a53af63db43e1946fd48e8459138272a132b202a8f21f81cf616fa12;
// music[1852] = 256'hcb13de0eb30aab0b76092d08ff08b609270b6709e008ea0b700c430c630e9211;
// music[1853] = 256'h0c12fe115d17781975166519201b8d19871dd01f2e2296285729fa298a2dcd2c;
// music[1854] = 256'h812c2d309f32f43091317c3391313b34fc349830c5334436fb37f639262f1724;
// music[1855] = 256'h0d24a62634269f25dc28b128d2276a281c2bbb3cb64985442943e044e344d147;
// music[1856] = 256'h024a414b1f4ba3495b498649f14725467c440042c042c84363447144a1371a28;
// music[1857] = 256'h1425f82487267f2bf8284923a9245e259f23a6229520cc234525bf22ce254c22;
// music[1858] = 256'hd91da5228b20001cef1d0b21c9219d1ec21ec71f9e1c971b6a1bf61c5f1d7118;
// music[1859] = 256'ha6170019aa18fb184d16e413ee12b5120814c9130e15b414580fab0c9f0e5d12;
// music[1860] = 256'ha813d413e512b60d260fba121d0ec00fd512a60e761037131413711370114a1c;
// music[1861] = 256'hda2980277529a02a3525b12be22e4929ac29142aa427252881296a28d7276227;
// music[1862] = 256'h27275d270b22f5206c213012fe049b056305510438067105c701c1012304ea02;
// music[1863] = 256'he2018e0336029101bc02bcfe45ff4303ecff8bfea3fec9fe4b030e0661074605;
// music[1864] = 256'h0803680482034005eb0758074a071f075808cf06af022d011a00840018049706;
// music[1865] = 256'hf4024b0137059402500093036b0420049d023703b90358fff2ff470395009afe;
// music[1866] = 256'h270321054e01170208033706d114381daf1c991d481d5420b722d920481f031e;
// music[1867] = 256'h65221c236a1ddd1cc41bf81da6215a1d491b4f1c2e1da3146d043304e0079404;
// music[1868] = 256'hf603b800700198022dfd10ffcd003bfd73005503effe08fdd8fe8fffc9010502;
// music[1869] = 256'h43ffa5ff6f007f01f903b106f806fb0186ffacff7c002902fafdd1fd1a0016fd;
// music[1870] = 256'h3a00ae015a00c80291fffefd140264043503cc00ba011b001cffad002000f604;
// music[1871] = 256'h2304ba018f0e0b15941378169317c718ac15af1388168214ea1d512b732a672e;
// music[1872] = 256'h84300e2b212f65319a2ec12e412f26318c2f382cd42c1c2cda2977295f287324;
// music[1873] = 256'h502483217e11c1047204160ab70c7d040dffd90045fe7efa5ff9a5f843f702f6;
// music[1874] = 256'hb1f62afb5efd94fa97fc5ffd74fa46fc23fac5f7a1f9adfafbfdcdfcabf7a5f7;
// music[1875] = 256'h3ef9a9f692f2cef3d8f0d5e994eb0cec8ae800e722e3dbe0b1e25be2eddf4ce0;
// music[1876] = 256'h5edf8edb10d9a6d551d787dad2d5ded2fcca52bec6bfdcc06cbdc1c12cc059be;
// music[1877] = 256'h6bc1d3bcf3c6c9db28db8ad7cedbb3db48dc28dcd7dbe8db5fdb9adf81dfbfdb;
// music[1878] = 256'h33ddd4dc80daebda17dd86dc9fdccfdeb0d0e5be1ebf7cbf43c07cc3f4bda1bd;
// music[1879] = 256'h23c043bdfebe58c1a2c2e4c5c6c574c354c504c7f4c365c69aca8cc61fc545c9;
// music[1880] = 256'h5ecb8ac81fc601c850c953cccfce82ce9fcf57ce7bcee7ce30ce72d1c4d011ce;
// music[1881] = 256'h35cc23cb2ccf2dcfe6ce50d186cf9cd21bd5f0d053d1dfd347d32ad2fdd2aed4;
// music[1882] = 256'h53d402d6b0d9a4d909d8ddd9c1dd3ddb77da28ea38f7f8f588f5ccf8c0fbf7fb;
// music[1883] = 256'h56fd17fed1f915fc67fd22fb29ff34fe33fb3afb37fc35ffacffd702e7fa10e8;
// music[1884] = 256'h25e45ae53ce5b6e7a7e68be4bbe177e2f4e4bae33be2cee0a3e0d0e2d2e5c0e4;
// music[1885] = 256'h64e259e237de4ddd99e0b7e398e69ee3d2e463e684e44ee9caead2ebc9eb5be7;
// music[1886] = 256'h7dea5ce93ce5aee6bce61ae737e497e47eeab8e71ee622ea7fe90ce844e7a9e4;
// music[1887] = 256'h54e440e51ce510e64ee764e842e82de6c3e7fdeb03ec6ce9bae9dae72ae572ef;
// music[1888] = 256'h72fe52055806a505ef082d08fe03b807100aa109150a6b08c4075b06dd04ef05;
// music[1889] = 256'ha8071d08fd06e509940994fa80eabfe812ec0fe921e714eaade9d3e922eeb2ec;
// music[1890] = 256'hefe90aed72ea72e89aedbdeb73e9a7eb2cec75ee2dec15e9eaeb14ece2eaebea;
// music[1891] = 256'h4cec59ed75ec1eef04efa7eb3ceb27e824e7a0e845e6fae617ea04ea05e9a2e7;
// music[1892] = 256'h56e65ee983ed2fed7deef7ed28e986e834e570e56feb94e920f21c0240049805;
// music[1893] = 256'hfd0581013c03ef063d04d6055c147e1e8720e4232d23fb228823bc215220e61c;
// music[1894] = 256'h041e982077203b23f221901d3c1ddd1d671b1b1d4322db1487037e057405d6ff;
// music[1895] = 256'h44fff0fd71ff6d01b6fdaafd4b007ffea2fff9ffb2fb80fc07ff3dfffffdbffb;
// music[1896] = 256'hdafd89ff48fe89fe1a0004011a001dffadffdb04d8067e008f000a018dfd88ff;
// music[1897] = 256'h7bff93000802a6fecdff5c0043fed2fdb3fe450106fd63f9a8fd88fc76fa4cfb;
// music[1898] = 256'h74f719faeefce0ef9ee80feb75e660e6dfe792e564e7c8e899f2d7fe89fe2802;
// music[1899] = 256'h8907db04ab030205a4069c07f5072b09f70a4d0a3f06f606430a2a0a22081604;
// music[1900] = 256'h7b053404ebf6ccefbeee1fe9bbe742ebe4ea91e9d1ec2aec81e849eadde95de6;
// music[1901] = 256'hb0e518e996ecb9e954eaecedf3eab4ea3dec1dec95ed91ecdcebd0eba6ea4cec;
// music[1902] = 256'haceddfed25ec61e8dbeae5ed9be9d1e743e88ee7e7e9e0e8dee6a4eaa3eb30ea;
// music[1903] = 256'hb1ea82eaa4eb3aede1ea52e988eb97ea23e9d4e90ce818eacaee2cf03fef99ed;
// music[1904] = 256'h09efcdec8aeebbfe7b09210aeb0a010e410fd80a280aca09630acd0d1d0ba30c;
// music[1905] = 256'h970cea09fd0ede0cad0ca40f1c0d740da20032f1cbf15cf0bded22ed2deb3cee;
// music[1906] = 256'ha5f0ebec75ea21ecd1eb84e939e96eead5eaf7eb72ee45ed5eed54ee2bea4feb;
// music[1907] = 256'h52ef0bf1cff16aedafec92ef4cee80efc9f284f23ef289f539f43cf1e7f219f0;
// music[1908] = 256'hf6ee19f1baed67ec6eed6cf089f20fed3bebbcee8eeedeecd0edb5f063ef61ec;
// music[1909] = 256'h2feef8eeb8ed73edcdea3ceb66ef1beef5f0aefd770627092109fd086d0e7011;
// music[1910] = 256'hb60c060b680e0110500e560c1a0ddf0e2e0f370e590e2d0f160e3d0fb708a9f6;
// music[1911] = 256'h45f1e6f386f0f3ef94ee63edb9ef91ee13ee3bf213f40df14bf1f9ee8ae8bdec;
// music[1912] = 256'h82f0b8f046f78bf98df938fb13fde7fd13f9a9f674f5eff1eff180f06ded1eed;
// music[1913] = 256'hd4f0f5f2b5efbeeeb1eef8eee8ef83edd0f050f655f5aaf48cf1b2f0f3fb5bff;
// music[1914] = 256'hf7f984ff6bfec3f82afeb5f8d3f84d0fce1847167c1a002067245f24cd224f2d;
// music[1915] = 256'he6403849fe4600491f4ac948f249454bf34a5147ed455a49d84c174b593eda36;
// music[1916] = 256'hbf3e9a41663fe947cc4c333dc02c592c102d5927d020041b8c19041894115a0e;
// music[1917] = 256'h0e0d9c090f0b910b0c0737051406140af10ac107370ab10a870d8d158d153317;
// music[1918] = 256'h961ad7187a1a741c4c1f972274223c25d9267e26042b432cd528402af42e4733;
// music[1919] = 256'hec3415323730b7311f352e36a837413d4c3c8f3cd93f853da13f4136f0251126;
// music[1920] = 256'hc626a529112b932642294c2c9a39e5478745df475e4aa248894a054a5749e348;
// music[1921] = 256'hed4863489145d145ad48f748b0434442c942ea400944cd3b352bd727c0287a28;
// music[1922] = 256'hae27c625f925012625269a25d5233b22ef20b9210423a022b123c8253124c123;
// music[1923] = 256'hc223451e8d1e0c226d1f881e69202f211120aa1f4a1ea11aed1baf19d516f51a;
// music[1924] = 256'h06183a16321af0187a184f16a41247144e13640f051174130311611297150a13;
// music[1925] = 256'h5712cb11cf0e830fc810da10f10f710f71124b14aa0f540cdf1a152eb62cac26;
// music[1926] = 256'h7328f028582b502d6b2c392c552a452a542a9b28852add28e523c4245d253023;
// music[1927] = 256'h3524fd20a1108204ce07df08360730072a023901770214014e02d5002901d502;
// music[1928] = 256'hadfee6feb3019c007a00bb004f00aa003c022c02b601e603520202ff89007c01;
// music[1929] = 256'h810174024d01230320073c04940376097d083a042e049d035403db033b038802;
// music[1930] = 256'h270240021e0369039001e5005f02cf00dcffac02fd012cffefff870051ff9e00;
// music[1931] = 256'h69023501b7089618f01d0f20e7223f1df61ef123ba20a621e322d92122221622;
// music[1932] = 256'h32236f2126209d208a200b20ba1bcf1a1913ed013e0041036fff1c0071ff38fc;
// music[1933] = 256'hecfd4502e6020a03210336fe8afeea029c025504ca0391005402c1030104d203;
// music[1934] = 256'hf0004d011c059f0698043f00affe25018e0199fe99fb7cfb5cfe590293048d03;
// music[1935] = 256'h2102e10221054403200044037e0370028d05df03570070fe52006703e300ec01;
// music[1936] = 256'h1203660740165c1959131d13a11341138612a51c582b3f2bca29e22bf5284e2a;
// music[1937] = 256'h382f9a2d982ac02be72b732bad2bc929092a792b812bd22a2328902968264115;
// music[1938] = 256'h470a7109d5086d0c100cf6038500b50070fe8dfce8fa87f910fad6f7e5f6b7fb;
// music[1939] = 256'h29fc1efad1fb26fd08ff930069006ffe88f9bff860fb02f84bf38af4cef5c0f3;
// music[1940] = 256'hbef262f152eef2eb24eb01ec19ebe2e8ade945e92ae613e55be247dd3eddffde;
// music[1941] = 256'h4cdd73dabdd915dcaddb48d933d9bfd4a2cabdc118bfb6c093c30cc4b9bfa9c6;
// music[1942] = 256'he2d522d75ed68ada0ad930d8bedb9ddcc2d9bcdbcdde77dba5da45db7bd9a6d8;
// music[1943] = 256'hb7d8cfda71d860d7d3db99cf9abde4bcf8bec7c0dbc4cdc12abef1bdb0be35c1;
// music[1944] = 256'h50c299c496c676c5f1c655c789c6a7c9d4c934c674c509c9f6cc6cca8bc791c9;
// music[1945] = 256'hc3c785c802cd47ca04cbfecd4acc3ace10cd89cafccb74ccf4cf93d10ad068cf;
// music[1946] = 256'h2ccd59cecdce8ecdebd083d17ccf0dd28ed402d361d389d5a1d43dd7a8d9fcd5;
// music[1947] = 256'h76d862dc0ed8c0d83edb7ddb61e971f7baf6b7f6d0f8eef799f936feb1fd1afa;
// music[1948] = 256'hcffcb7fcc9f99bfb9efb2bfc0efb65fafbfcaffa04fc8bf73be8aee4cae512e5;
// music[1949] = 256'hc6e646e57ae3eddfc3dd62e058e145e38ae4a9e252e3b1e306e09dde0ce3dae4;
// music[1950] = 256'hc8e2e4e4b2e8c6e9f2e9c2e86ce6b3e640e70fe5a2e5eae632e597e551e7eee7;
// music[1951] = 256'h00e67be4d2e62be592e4c4e9d4e7f3e4bae9c7ebc7e960e9c2e766e681ea27eb;
// music[1952] = 256'hcfe68ce785e8c6e9eeeb9ae7d2e5b9e904eb59eb07eaebe55deb01fddf04a401;
// music[1953] = 256'h7a0416049fffdd0304075b04bd05f2082d0835079b06b90502077605a6028203;
// music[1954] = 256'h0206be0572f759e721e90deb30e774ea39ec73e930ea48e972e636eae3eb8fe7;
// music[1955] = 256'hfce905ec45e7fee6eae796e727ecd0eec0ec86ecadec57eb43ebafec15ee61ed;
// music[1956] = 256'h03ebe8e99ae888e6c6e61ee762e68ee832ec84ed64eb3ce8eee8d9eb2ced4ced;
// music[1957] = 256'ha6ed8eec4fea01edb1ee63edbcef96ee2eef3ff240ef90f4d4fe760467061d02;
// music[1958] = 256'he5026c020902941473215d1e9f1d761c8b1b831dd91e561e6b1d9e1fef206121;
// music[1959] = 256'h68209a1ada17f8170218a119191a411a751345079002550204046e05fe046c03;
// music[1960] = 256'h3afdb9fda401fbffa70172fff3fca201d801e50091ff13fd3cfeddfef5feabff;
// music[1961] = 256'hd0ffb2ff2b017b0226ff0dfcabfa5dfb05fec0fc42fb31fbb8fcb500cbffb1fd;
// music[1962] = 256'h69007f01a7fdfffa9bfdd7ff7afe1bfe99ff2bfe0efc72fd85fdbcfbc4fb15fc;
// music[1963] = 256'heffc56fdf8f56debebea7fec4eec91ec02e74aee38001002c3006e023700f601;
// music[1964] = 256'haa04b705e30661065b0537058704c1015f021b043d021f017d0010045203cff1;
// music[1965] = 256'h07e769ea7ce952e995ea74e7eee63ee75be60de7ffe6dee68ae798e817ea86e9;
// music[1966] = 256'hcfe8b4e96ae840e820eb36eab9e83cea5bea54ead7ea81eabdeaedebf0ea7ce8;
// music[1967] = 256'h8bea90ea4de7c6e807ea84ea76ebe4ebb3ec85e931e933eca0eb23ecf6ecf8ec;
// music[1968] = 256'hbdebf0e999eb77ebe2e9cee920eaa7ed6df1b7f088ef97f03bf033ef53ee46f3;
// music[1969] = 256'hda02e9081e055508e707c7055f09da0a310b640b070ce20b5d08f20654087508;
// music[1970] = 256'hb006870666064b06250a9e0215f10bee62f099edbced2fedf4ec69eda7ebbdec;
// music[1971] = 256'hacec37eb0aeb47e926eb8dec71ebfced9cec15eb6eee74eedeee82efcfed06ee;
// music[1972] = 256'hb3ec5dec75ee7ded07ed0bed20edb1efb8ee52ece3ec6aec4eec20ec77eb33ed;
// music[1973] = 256'hbdec5fec52f0c6f186f1eef03feef2ee6df04df09af06cef00f14af3daf293f3;
// music[1974] = 256'h88f407f519f362f200f2f5efb6fcc50a4108ee064407b1074f0bdd0a8e0b8d0d;
// music[1975] = 256'hd30c770b8c091f09a309020abb083609650bde081b0a5d0853f7deed63f103f1;
// music[1976] = 256'hebefa9ef15ee66eeb6edcaec72ee0bf074f0bcf103f360ee23e9c8eb3befcbf2;
// music[1977] = 256'h33f8c8f846f8fef9cbf846f7aff79df5fef259f294f1aff04cee79ed7ceebdec;
// music[1978] = 256'h08ecd2ec74ecd4ecf5efb2f2ccefb7ee59f11bf3a1f5d4f9240208058900c0ff;
// music[1979] = 256'hb6fdbafdea00f3ff89ff6a039010161e3a1f7f1f78225d24912e013f4546ec44;
// music[1980] = 256'h0f439e4209462249ca49ba4a204a3b477d453548a54aa248f53c64310a3ae83f;
// music[1981] = 256'h8e3e17457d3bf12d3b2ddb28c726ba24eb1efe1a7916bf13cb10280c9e093b09;
// music[1982] = 256'h5f088505fe055e07f2053006ac08b70b730e400f5e0e3e1041134f12cc139e17;
// music[1983] = 256'h69174f17561a7c1d3f1fbb20a0226d24f625ab27cc29bb2bf42c9f2c822da22e;
// music[1984] = 256'h1e2e0c31063382333b36b135d0368c39e539dc3b223de83f363dd930a82a212b;
// music[1985] = 256'h7a2cab2a442aec3836453245f14491423a43e2451f4491449a4469431544b945;
// music[1986] = 256'h4147dd45244561431542f8439c410942c73ecc2ec328f42b382a6f281e270b25;
// music[1987] = 256'h4d23d7236424842105200a21692221229720e220c72096200520201f0321e920;
// music[1988] = 256'hfe1ebf1e341db61b5d1a1d19dc1966193f186d182d18c717a71649159a164b18;
// music[1989] = 256'h0a17fa157a16a314a2121213da120d146516a6164016d514e314e9155d148e13;
// music[1990] = 256'h7712aa120214e7117b133614cf108e1105104116dd263b298d25e42676258925;
// music[1991] = 256'hf426b725cd22a4225e240623cd246225012295214020ea20672132218721e613;
// music[1992] = 256'hb20777097708900772075205af0451038f0460052603970330043a034d039103;
// music[1993] = 256'h5d027d03dd0428029203c606130529047004a804c4036d02d3035d03b9012402;
// music[1994] = 256'h0202f801920132015f028d0264027e02c40002ffa9fd02fc20fe33015200e900;
// music[1995] = 256'hd802fe02d905b008bd076f0717078e054b06b9068906210798059e051505b006;
// music[1996] = 256'h6515af1e941a971b8c1ecd1e6b1d7b197919691cb91dc31cf01c181e351c6f1c;
// music[1997] = 256'hf81c691cbb1b0e1ac91d97164b03df00270462001500fbffa7fef7fdd0fea400;
// music[1998] = 256'hb2ffbaff560055ff66ff0bff26ffb0000701cc00c2007801d6020b025700ab00;
// music[1999] = 256'ha702fa04e8042f02a5ff48ff5d001e00c6ff3b0061007200ceff8400c0013f01;
// music[2000] = 256'h08020f031503b5035704300481047906e9070d081307b706cb07b006a8054f03;
// music[2001] = 256'h6c086c19001b3f154f177f12f11a332c022c5b2bd42c662b4b2ab8266c270228;
// music[2002] = 256'hfb26ed29d52acf2a162a6e2840285727fc255b24d7264a25c914fb099b095903;
// music[2003] = 256'h0801d8078409b0055b0357ff92fa80faa9fa6ef81cf83ff924f9f0f83cf9e4f8;
// music[2004] = 256'hbef956fb47fda5fe1dfc7afba3fc3ef9e9f66bf786f717f51bf26df201f14def;
// music[2005] = 256'ha4ef13eec9ed16ede5eae2e9e7e7ace46ce0bbdd48de91dea5de33e11fe262de;
// music[2006] = 256'hbfdd47de8cdcbfddbfdbb2d92dd9bccec2c3aac288c3c3be68c0c5d13fdbffd8;
// music[2007] = 256'h7fdab1d966d656d5c7d4b9d44bd52ed6aad603d887d681d5d4d7cfd5c2d695d8;
// music[2008] = 256'h19d77dda28d227c288c14ac2e0bd09bff0c0fcbfa7c065c1e5c0e1c104c2e8c1;
// music[2009] = 256'hacc3b5c3c0c3b7c5a2c62fc6a7c6c2c6ddc609cac6cad9c87ac9d2c84ac8a3c9;
// music[2010] = 256'h0aca9ec9b1c9f6ca01cbd4cb99cdfccc24ce3ecf72ce37cfc9cff2cfbfd0d3d1;
// music[2011] = 256'h6ad272d4d0d713d8b5d84edae0d99fdaccdb9cdbdfda9adba6dccadc0cdd45db;
// music[2012] = 256'h72dcb7dd98dc89e8dcf4d4f40af7e8f63cf3d5f3b4f2c9f02ff1a7f2e2f3ccf3;
// music[2013] = 256'h44f41ef5ddf5f9f469f4faf525f63af89bf57fe7e9de98df9cdffbdf5ae002e0;
// music[2014] = 256'hb2e0bae165e1e2e0bbe275e3fbe2dbe30ce3f3e2e4e3e1e1a4e18ce32fe30de4;
// music[2015] = 256'h44e6f5e6ace7c9e746e729e75be6cce5bfe59de504e67de687e69ee615e754e7;
// music[2016] = 256'h7fe7b1e7dbe7cfe84fe942e819e632e62be921eae1ea6ced32ef71ef30eee1ee;
// music[2017] = 256'h00efcced1befddeef9ee58ef64ee14ef2fec3df055ffc30584041203a301d102;
// music[2018] = 256'h66026b00a2ff79ffc5ff64ff7dff78ff79ffcbffb8ff4901b600aa00e3022df9;
// music[2019] = 256'hcaea1de8f5e8eee7cee724e861e80ee8bce89de9bce93aea34ea29ea4cea3cea;
// music[2020] = 256'h40ea3fea48ea2fea80eafeea49ebe6eb86ecbcecdeeb5aebb1eb94eba1ebc5eb;
// music[2021] = 256'h3deb37eaa6e96ce918e933e9ace942ebd3ebcdebeaec39ecddecd0ed57ec60ed;
// music[2022] = 256'habee2bef01f13ff28ef2e3f2e2f2a8f196f22cf12ef295008e08c106da065e06;
// music[2023] = 256'h1e13b020421d7c1b891c1a1b1b1b181ac0180b1805194019df188c190a196719;
// music[2024] = 256'h5e18d8172719cd17c4193215770413fea2006dff92ff3400cbff8b002f00bbff;
// music[2025] = 256'h1f00faff12002a00d1ffbdffddffb6ff33ffbbfe97fe36ff68ff41fec7fec700;
// music[2026] = 256'hf1007a0046008fff38ff1affc3fec4fe9bfe52fe98fea4fed5fd51fcbffbaafc;
// music[2027] = 256'h95fcadfcc5fe2f0049ffd6fd5efe0affd3feb800b801c000d600b200bb00f800;
// music[2028] = 256'h670100fc01ee4eea3ded5de952f2560118023a0150021902ef02c00256026a00;
// music[2029] = 256'h6cffb20084008f001d002800b9008800b501a600df0141024cf4b9e8f3e909ea;
// music[2030] = 256'h35e952e961e891e87ee82ce803e8b2e725e8abe863e94beaa2eaa6eae7ea65eb;
// music[2031] = 256'hefebe0ecf7ec38ec48ec97ecb7ed9feeaaed29ed4aed18ed24ed40ed23edabec;
// music[2032] = 256'h72ec87ecb0ecd3ec8cecf8ece0ecbbec25ef76f0f3f00df259f062eff8ef40f0;
// music[2033] = 256'h66f2b8f290f159f1c6f015f14bf0feef8ef06defa6f07cf071f3a900b0074106;
// music[2034] = 256'hb5062c0675059c0593052e05e903930460054a059a055905db053f06e7060807;
// music[2035] = 256'hfb05fa06240005f2feed6def89eee3ee20efcbef00f0b5eed7eed7ee7ceea8ee;
// music[2036] = 256'h14eebfedc2eda4ed04eea5ed03ed67ed4cecf6eaffeb8fecf0ec54ee47ef4cef;
// music[2037] = 256'h79eea6eec3ee8aeea6ef8aefceeea0ee1aee4eee3aee52ee24ef4cf03ff227f3;
// music[2038] = 256'hdff28cf2adf1c5f084f05af18df389f58bf55cf568f5e7f499f487f49ff470f3;
// music[2039] = 256'h2ff445f62ef545fc45080e0acb08e308780844089f07aa07df05b70450051205;
// music[2040] = 256'hd305eb05d306f90696064408690537056405a5f8c1ef44f12ef1fbf0abf1e8f1;
// music[2041] = 256'hf9f13cf112f1faf0b9f072f1faf27af543f58aeef6ea6aef2df2cbf344f759f8;
// music[2042] = 256'h01f984f954f85ef7dbf6d6f62df6a8f49ff311f2bcf0fdefbeee7bee38eff1ef;
// music[2043] = 256'hbaf01af1eaf132f4b3f6a3f7a8f74ff728f7b5fcd403e50196ff3a02aa00aefe;
// music[2044] = 256'hc2fff800ef048707b9088a116d1f3c278225f528803832414d40fc40ae41d841;
// music[2045] = 256'hab4190412941613fd93fd93f5b3f30418b44a44291340b2fa2357836f73a5138;
// music[2046] = 256'h662a3729ba296b256a23481f891c56191b15bc12b60fd40d5d0bd5081008a107;
// music[2047] = 256'hd0072d070e07b907f6077b09d70a300cce0dac0e1710671297156b189519601a;
// music[2048] = 256'hac1b121da21e5820ba201821fc22462404266329c22b592dd02e722f84307531;
// music[2049] = 256'h2232e23288322534de36c93759388837d537ac388e39033a74314f2b0f2cda29;
// music[2050] = 256'hcb333a41d840c040ce414a41e44147413841024010402e41f1402d4225425442;
// music[2051] = 256'hd641b33fbc3f693e9d3f6a3d7c2f3928cd29c5284828c627c326a326b1254e25;
// music[2052] = 256'h1425fd230f236d22d0217f214c21cf208120f41ffb1e281f6b1f691e1c1e9f1e;
// music[2053] = 256'h6e1e201eaa1d071e1d1fc61d501c241c141b861aae19e318281908180318f019;
// music[2054] = 256'h241a43191c19ec18c618c7191d1ada18c9178f167315fa14dd1487141114d713;
// music[2055] = 256'h4e139d146a1542147f13720f18136b21aa25672337245123aa222a2278215c20;
// music[2056] = 256'hf91ec71fa01f371f4e1f8a1f6e1f7b1d991e971ec71d921f92150209b608f008;
// music[2057] = 256'h3c08fe088f0820094009ab085c081c088107e6067e072f07ca06c20677054605;
// music[2058] = 256'h4d059b047a040804fb03e403e802df0156019201220230039103d602bf026902;
// music[2059] = 256'hd901bf01e6017c029f02b303ee04c90465056d05880582057503b00335042104;
// music[2060] = 256'h45069e057d049805f9045604de0480065607a9064b07ae041404c70fcc193d19;
// music[2061] = 256'hfe18cd192d19e318b017df1665162d160d173917b0174d17ac1521151016a616;
// music[2062] = 256'hc615ac171e133f04b0ff29020b0148019a0042019e02fc01130355037003ad03;
// music[2063] = 256'h5f03b0035503870390037503e203da031304bc031704cd03f601a2022f05ec05;
// music[2064] = 256'hb80362029c0270022f02c8002801a5025a022402fb01e9035905d404c5056f06;
// music[2065] = 256'h1c07fc0627068d06d7059c059c0628081d08cd05970533064f065e07a5083f0c;
// music[2066] = 256'h6c1391160b1277161223d5244c22e422ee224223d122f621aa20bd2081215021;
// music[2067] = 256'h7122c620a41fb920231f6b1f6d1ef11d021ea5119105c4044103240042021b08;
// music[2068] = 256'h6d07ee0142004dfd3ffa33f92df7a7f769f82df8b5f831f95cfadcfa9afb9bfc;
// music[2069] = 256'h51fc99fc8bfc37fc8cfb44fa8cf98df8b9f7f8f6a1f671f6cbf3b6f0aaee1ced;
// music[2070] = 256'h55ec72ec2dec21ea64e828e7e8e540e5bde331e2a6e0badf8ae012e088dd97db;
// music[2071] = 256'h4cda98d997db0fdbefd85eda88d2a9c509c275c423d0bdd963d722d790d700d6;
// music[2072] = 256'hbad633d658d47dd3e9d459d547d42dd301d223d387d35fd486d53bd435d6d0d0;
// music[2073] = 256'hf7c2d3bfc4c172c0f8c051c12dc128c2c5c246c3f4c35ac4ecc49ac553c6e9c6;
// music[2074] = 256'hd7c68ec78fc8c5c84fc95bc9a6c99fcac7ca99cbfacce4cd77ce61cfb7d1c7d2;
// music[2075] = 256'hebd178d2bad392d39bd239d2d9d286d411d60bd6add5a9d5dcd5fad6c7d864da;
// music[2076] = 256'h3ddbd3db93dcb9ddd3dd14dd4bdf1ee01ede52de84dee5de89de12de1bdfa2dd;
// music[2077] = 256'hafe59df339f51ef5dbf641f654f7f7f53af404f498f431f584f3d5f35df4a7f4;
// music[2078] = 256'hc3f571f506f713f7c0f72df7cdea49e2e8e30ce3bbe238e329e279e21ee3e1e3;
// music[2079] = 256'hf4e380e3bde38ae378e342e4c9e417e56de541e548e5a8e5d5e512e751e838e8;
// music[2080] = 256'h58e8cfe841e9e2e91aea18e983e71de7dce774e91beb59eb13ebffebc4edb5ed;
// music[2081] = 256'h50ed14ee64edaaed44ee94ec9eec70ed7bee8ff0e0ef2def09f15cf1bbf074f0;
// music[2082] = 256'h1cef91ef12f059eef6ee5eedadef42fe6305e202aa03a3037e0333036f014b01;
// music[2083] = 256'h4701300030fea3fe03ffd1fde8fe86fe96ff1a016600cc024afb2ced84ebf4ec;
// music[2084] = 256'habeb5cec09ec72eb4feb67eb13ec1beceeebd1eb7ceb37ebd7ea57eaede9e8e9;
// music[2085] = 256'h7aeaa7ea21ea6bea0aeb39eb99eb4feb90eab6eab8ea4dea13eaf8e989ea52eb;
// music[2086] = 256'he8ece5ee94ee10efc6f017f0ddefdeef5aefabef3aefeeef19f0edefddf234f3;
// music[2087] = 256'h83f2caf433f648f689f56cf5def3baf2a7f30df1e6f7b40296013d0bec18d217;
// music[2088] = 256'hd917261872175c18df1522165a16de141f150415181545143514e813d813c915;
// music[2089] = 256'h7814261682140d069dfed200bcff43ff53ff13feb4fec9fe11fecafe8ffe2bfe;
// music[2090] = 256'ha0fe62febdfe6eff69ffe4fe7bfef0fecafeb9fd62fd01feeefd43fedcfeadfd;
// music[2091] = 256'h93fd2afd11fcb2fc79fc0ffdfdfc7afb32fc1efd45fe5afec7fd4bfedcfdcbfd;
// music[2092] = 256'h72fd70fd9dfd64fc10fda2fd58fe6a008200ceff6f009800050097002dfff0fd;
// music[2093] = 256'h72fc72f2b2ec1cee00edbeed60edd2ed2eeeaeee1cfd30086b05b6050307de05;
// music[2094] = 256'hce059f05fb05a406c506b606f8060b07e706b006990643066e06fe06a705a907;
// music[2095] = 256'h2b0513f48cea60ed59ecfbeb01ed90ec0eed98ec87ecb6ec67ec79ec16ecbeec;
// music[2096] = 256'h58ed3bed18ee20eee6ed5aee2dee8aee43efbcef90f00af17df126f1f9ed7fec;
// music[2097] = 256'h13f29ff7d3f6b4f44bf4f9f421f5b1f234f022f35bfb8ffebcfb7ff900f5eaef;
// music[2098] = 256'h85ec83e850e704ec2af3c0f1efe314d504d4d5dfeee5ade0f8d705db13efbcfc;
// music[2099] = 256'h32fba2f5cbf8f9038d00e6f99b03d50f6313fa0553e91ed100d465f3cf0e7218;
// music[2100] = 256'h2a1b8919e3160116d912a70e7b0e1910df1103145c1b4126381799fabcf90c07;
// music[2101] = 256'h6d116c12d102c5f9f702a3116617060988ed4fd8a7d583e62204441fb528fc1c;
// music[2102] = 256'ha205d2f2feee72ff4218e21f251273fd0ef2a2f253f4e7f235f0f2f0aaf6a604;
// music[2103] = 256'h2e180a1a4f0fcf0e4e0e8d06c4fb09ee1eec39ffde17fb211a1a910f59096d01;
// music[2104] = 256'h79fbbafb32002608db10fd16cf14b50421f162eb8af011f839047710121dea2a;
// music[2105] = 256'h3e324438b33bec3e3f5267680a6d4560594fdd46203e902f901d1f0522ebd5db;
// music[2106] = 256'he8e3c1ef69e851ef620e7820d01f100c65eb53e06ee63ee5dde42eee01fe7508;
// music[2107] = 256'haa097a0f6118941e502b6a3dd9453041b63f4c4c0e5ee4653661ab5979598c65;
// music[2108] = 256'h7d64924abd41d24c7b494a3b13328632cb368a4384571c52a1342627ab3b4857;
// music[2109] = 256'hf55517493247ae441442864c7763926b24543d3557295c2e752f182b0029e026;
// music[2110] = 256'h4727e425782c0442ef4f65557d5a4054b73be61b070830fed9fec1071efd84e9;
// music[2111] = 256'h97f6a91ec837f831382cea38f335311ae10b3617b33667517846dc359840ee4e;
// music[2112] = 256'h1f49823bb13f48402e2cd61efb1d69237826151b910caf11ad2663261717121f;
// music[2113] = 256'he12e2b274711790fc81f3628b829c824ff1571062e08de1c80252f17b4ff35f1;
// music[2114] = 256'h7af4ccfdbc053b089a0cd1175e198512e506d8fbd3052e1caa26272747189af0;
// music[2115] = 256'h89d009c867cd88ea5b0531fedbe1f1cf8ddceaee2af85b00b3062412811d8325;
// music[2116] = 256'h0720750061e298d332d577e6a4e729d845dc58eea1f7f001570569f462e6f8e0;
// music[2117] = 256'h67e07beae400ef19f8150efa55e5bbdaf0deeef28f130f34e239742746088fee;
// music[2118] = 256'h20fc751ddd295327a71fe51b44268e30673b743fd52be11dfd221e3121449b39;
// music[2119] = 256'h380cafe804e9d307fd272032182ff2265f1f9d28a42bd109a3e449dfd9f68a18;
// music[2120] = 256'h1c27ed1e6f121d075bf544e2f0e597facb07e20dfa0c8608f009d00525fda500;
// music[2121] = 256'h5605150538ffd3e3ffcd8cd7a2e049de47dce2d8c2d863ddc4e120eff9025dfd;
// music[2122] = 256'h7ce410da69da06ea9b04c307b9fa19f5ddf368f31dfb0a08ab0eee1455198017;
// music[2123] = 256'h1815710b8d0834198324f01ce20f340511fff40e0f273d1be0f9c9e86cf3a711;
// music[2124] = 256'h17207c18051c642af52bc222b81983182e292c3af435632924253924e5215828;
// music[2125] = 256'h9c2a9f230d308444de466f338e173f10371b2d2c4a338d28a02cc341694e834c;
// music[2126] = 256'ha14cf1596658654f304b2634b72293273c21940230edb3fe9c140d174318bb1b;
// music[2127] = 256'h68215b1e430f2a0c401458213a2fbe29c51ee41a570f6606fcfb08e905eac703;
// music[2128] = 256'h9c126703ee04ef288a3aba355a27691a74263f337730a823df1c2620ff05c4e2;
// music[2129] = 256'h3ddeb8f0f90bf60748e85fd3d9d0afe57bf3daea93ec3af3d5eedde6cae3fde5;
// music[2130] = 256'h4ce3dedbc8d2e1c655c124c1e1bf22bd5dbaa5bfeabe36ad72a351a9beba08cc;
// music[2131] = 256'h0ec9ccbf3bbfc6c5decac9c6f5be90aa4a9a56a2c1a9b2aa68a6eea249a8d0a7;
// music[2132] = 256'hbaaddcb7e2bd24cd62ce26c25bbdfdc01dd20dd8f4cbd6c062b3d8b2abb7acac;
// music[2133] = 256'h78a916ae0eacb4a78da1c9a952bbf5bf86b631a391af29e2eff92efc3f074f00;
// music[2134] = 256'h6fe0c8c565cf7af5f61248200827d622bb11ee05640aef0ebb03dcf4cffc581c;
// music[2135] = 256'h5a3c7941172b611b7215b31253196e126000bfffc412a2299932cc30a2301837;
// music[2136] = 256'h253e033df239402c6f162b109f18532d0e41963b1d2b40293b2eb125db20f534;
// music[2137] = 256'h81481d454a3e30455548fc3f1a3a253793310c26ea25143dee4d5a4cc6475e4a;
// music[2138] = 256'h234db53df527011efa1a0721fe33f54888526c511c4fa84c9a3d092c0531dd3a;
// music[2139] = 256'h053a5e375c3164318c38204775612d6c645b4e4bfd54596d6d793c75ed620750;
// music[2140] = 256'h77520d68bc77606ae84a4a387544a4615470de67f54d953f114f25555e446830;
// music[2141] = 256'h221ce8139c1e52300f3ff43b5a21b20d631579223a27b7285f2e5230971bf202;
// music[2142] = 256'hd7fc25faa3ef94e790eaa2ecade9d6e987eab0e9c6e7d7eb15f043e592dc9ce0;
// music[2143] = 256'h25e66fe2bfd4a3d060d133cd03ce25cb4ec866c9f9c2eebf32c25dbf06b893b3;
// music[2144] = 256'hcfb444b162a9b5a461b02ecc81d130bd7ca87a9f07b153c495c32ec089becfbd;
// music[2145] = 256'ha5bacfbd60d199dc68da27daecd95ed962da2bda32d999db29de92dbc5d95edc;
// music[2146] = 256'hd2dea6dd8cd9b1d443d60ddc68da2fd8bdd338c676be94bf41bfffb07c9edd9e;
// music[2147] = 256'h4da34aa3cfa5f1a3119b13961fad24cac6c8d3c3b9c74ec90dcacac89dc715c3;
// music[2148] = 256'ha4c1cac6a2c80cce77d491d787d782cf77cee2d4a8d2a1cf97d496d8d9d768db;
// music[2149] = 256'hf6def6daa6d8dadb4ce1d0dd61c610b37ebfdcd737e3b4e4bce081dc2cd41ac1;
// music[2150] = 256'h79b514bac8cde7e79cee32e756e5dbe8d0e9d7e146e005e7f2e8f7f4f4065205;
// music[2151] = 256'h7dfb05fe8f072d0efd0f9e10b314c1187f15d209c204630d870fd60ce50daf01;
// music[2152] = 256'h71f17bec45ecf7ee4aea7de86cfefd0726ed6dcfa0c6d0d215e05de49ff0b1fd;
// music[2153] = 256'h5202d004a602dc022308870b360894064f1713220418ee15fe1cee23ff297b27;
// music[2154] = 256'h4323a425f8298e2b8d2af52c0837af3a2a224b02e202fb17c128143389296512;
// music[2155] = 256'h5e0aa50e1310811250232a39633455169efee605c1222132d230cb2f1f32fd32;
// music[2156] = 256'he02ef52dfb2e462ef92f0432c631442b4f302d4d275ec4555451075a155d8b5b;
// music[2157] = 256'hbe5c9c4c69370a382c3b0636cf34423a91418344894bc35eb5634d4dc73fd73d;
// music[2158] = 256'h4131ae2a0b2c4a2985254228be3cd14d6a4f5855d45795563c593253f8499848;
// music[2159] = 256'h704a6b46bf426147614665426e439644b448bc45eb360826dc20d83792514452;
// music[2160] = 256'h154903474f4a233df524f12034236b1b6b1f91344a4478448941b644cb404629;
// music[2161] = 256'h6614f91b9a34663e873590330a340c2d5e2ec9342a366731ad2f3231a828d723;
// music[2162] = 256'h2f270a2e7131bf180807e01659215f1d9c1b9b2ecc4da351cd39d921b71fb733;
// music[2163] = 256'h8c47d045542ba019f622b533234238413f2a7817fd16d511e300f3027c16d71e;
// music[2164] = 256'hbf220f299527c221a51a29142116bf1b2b1c28192c19e51ad70a9fee52e8acf5;
// music[2165] = 256'h0e077b12d4036cea46e207e2a9de68df04e348e20ae369e2e2dafad7feda9fdd;
// music[2166] = 256'h05dc53d513d1e4d81ef1b2fc10e882cde7c119d28fe931e7ffdfe0dcc1d9d2de;
// music[2167] = 256'h00e149e012d926cf40d2a5c58aabaaa982ae04a829a4e7a51fa3099f70a91bb8;
// music[2168] = 256'h64c587d68bd587cbe3cd9cd2a4da58dadfcea7cd50d15dd3feca17b3a0a360a2;
// music[2169] = 256'h32a071998a9d5aa931a8c5b122c2d0b00c9d0ca0a8a2e7a514a978a26b946888;
// music[2170] = 256'h0388099047a08da649985b948592d48876883c8440854a9162984d9f239fbb98;
// music[2171] = 256'hf0958f97d89a699aa69ba793e086378730893694429d6590a68b5a95a592b186;
// music[2172] = 256'h34841586688ded9d739c1e92619004891286198857863788ed868b896d973996;
// music[2173] = 256'ha9865e85b58755857c865084e68c839f3ba4d9a16fa0d4a698b649c09fbcfeab;
// music[2174] = 256'h24a081a357a564a137a61bc0fad710cc61b1baaaedaf61acbaaa5dbfecdbc6e4;
// music[2175] = 256'hc2d4dbc15dbf42c600d4addaddc6e6b46db55ab75eb613ba7ecfa4e4c7dffecc;
// music[2176] = 256'h32bc37c227df0ef039eed9eecef7d0f3c1db2dcce7d2ece7aafc41fc16e9d5dd;
// music[2177] = 256'hbcdf70e0e3e20cf154076110d2009af1a8f2def616f352ee5df37df8a3f8c9fb;
// music[2178] = 256'h78fe7e019f127d2af22d471cdb086d04060c670988058105deff810716219e3c;
// music[2179] = 256'h06410927c50ebc05a80cf4169815151db7281a31c74c0d620356e442e63aa33c;
// music[2180] = 256'h3839bd2fa643d464e76e9270197108716c6be162d965cd58b5442f45f33b7b29;
// music[2181] = 256'h8a2d11457c589a5c575b145d975db95232448f3fd73fba3b813c0452f966ab67;
// music[2182] = 256'hdb67c46b605f0d43fb3a7b4a464b79421d4f216b9f75cb663f508047365cf773;
// music[2183] = 256'ha1785871bf68e06a78634e50754c07582d6a036eca5bca483d453e557b6a366e;
// music[2184] = 256'h09590d4797499456a165545e7846263b8843b45fd86e895f29442133403d3253;
// music[2185] = 256'h1864b15b0f42b5460c54634e9449f648be4786451251d4690d6fa15dd94c6646;
// music[2186] = 256'hcf415d3e1c410f402b3c763d8e3e81407f448b3a6324a51d0122de1ef41c561f;
// music[2187] = 256'h3921371de1115a0b3f0d11186e209b1a851476098efeba03f4070a18e234a836;
// music[2188] = 256'h6c282d2a4f3358279f0dc906160b7207f000bd09b31e9129f72d632ba122cc22;
// music[2189] = 256'he122f91f2d1e561acb12250d30146b19dc18191d12180f0b7f043406850bb30e;
// music[2190] = 256'h160c65021cfdd401e00a090fbefea9e0c3ceacd6b5edc6f952ec50d8eedf4ffa;
// music[2191] = 256'h8f0a090959f2e1d76ad661ed7a017902dcfdbdfc80fd90fbb7f53af4b9f97ffe;
// music[2192] = 256'h2af9acf329f49fee3fe868e1b4db45daacd35cce0fca07c619c8a5cc6dd68bcd;
// music[2193] = 256'h59ac579eaca451a811ac32aae99f74997e983f9ad29e47a7e0afcbad1eaa5ea6;
// music[2194] = 256'h75a0c5ae37c241c64ac9b9c835c429c12ebe09c0d0c1c4bec0bf5cc38dc124c0;
// music[2195] = 256'h6fbf3bbe8dbf20bc02bb6bbd05bdf6bfc3b5ee989b86b995a9b3cdb95cb376b4;
// music[2196] = 256'h3fb63cbae5b9eeb455b6d6b67eb28eb583bbcbbbacba29afd3a9b3c074d41cdb;
// music[2197] = 256'hc0e0adde7bd61ad010d61ce3d7e38dde9ddec7db38d74cdb89e1e3e5fce15cda;
// music[2198] = 256'h21d7a3c0f7a682a364a5c0aa40a788a7bfbd21cbefccf2c679c1f3c9facc7bcd;
// music[2199] = 256'h5fcccfc877c8acbaebb00cb648b5a0afaab1e6c57cd92adb26db79db8fdab3d9;
// music[2200] = 256'h96d612d6d0d409d716e0c3df76da75dabadba6df4dda95c73fc03bcfe1e545ea;
// music[2201] = 256'hc8da21cad8bf57c979deb0e606e694e431e985effceefae92cd79ac231c5d2db;
// music[2202] = 256'hb3f211f331e1fdcbffc65ce52b03d9085c0d73113612a6100d0bbc0810081c0b;
// music[2203] = 256'hb4115815471cd2180803bff82ffaeaf864fb16fc57fb55fa8ef08ee5cde258f0;
// music[2204] = 256'h6f05750f82112613aa1369041def43ed84ec9ce70de7d4eb80f9e3fd9dfcd7f4;
// music[2205] = 256'ha1ebc8011a182d1dc7203b189514c31b89259f2a03247f1f211273fc81f78004;
// music[2206] = 256'h9718f7208622ab28c72b372781212d21ec139bfe17fe2511c8290a29e90e31fe;
// music[2207] = 256'h52009611ca1ec420b9247029de2e772e42248b18400bc3fd04fc5e0d6c256f2f;
// music[2208] = 256'h1f2ed835de382f2fcc3587398427581c871bf1168b10c720573ca4424e44f046;
// music[2209] = 256'h9744fb398323211af71aa21c2d23161f6c0f3a07370d120dbe0a231a18244522;
// music[2210] = 256'h64222129252f0920990700fbaffa1700040a93214232582ddd28ac293920790f;
// music[2211] = 256'h8a0c73170427213278251911090d611a153217377223750dd4059b1b3f37613a;
// music[2212] = 256'h1e320c2b9d27662a7232f1372b28530dc108ad1f8937a13198152404eb09f11c;
// music[2213] = 256'h3a268c20b016ed0fd313f41f262ee029730d5804870bd2016effd80c88140917;
// music[2214] = 256'h9918121c8d1b8f12ec0e14119013cd12ce0e761e4c377e39903205333931d31e;
// music[2215] = 256'h5b08fa0ab718261295fdbef4f3f5f5f3bcf69ef95bf746f8dff61af42af5cdf2;
// music[2216] = 256'h33ec92ebb5f3f7027414d0150f114b14bb138514ce15ee155f183715ef137110;
// music[2217] = 256'h870f06173c0bd0f335ee65ffb5173219350314edc7ec1905691ab81fa4202b1a;
// music[2218] = 256'ha91044167c1e301dcd1984148d17ad220c291027c6215a21a6167e01edfc830f;
// music[2219] = 256'h1028702a871fa9193712f5126a19d31fa42d143be33cae26840cde0cce134f12;
// music[2220] = 256'h8110800c9109560d6413c113b5138424a8370936372fa42add270930c530481d;
// music[2221] = 256'hee0dc812311896169e1be517110372f33bf449f896f4a8fd6413961ae1157813;
// music[2222] = 256'h541454134b1487130106ddf9cafcf80c7615ce099a009a06b2145e1d461dff13;
// music[2223] = 256'ha9f5cbdbeee4db028b14810ffb075107a509490ab3063e047104a605a2f6b0df;
// music[2224] = 256'hcadb4ce590f4c5f9deeb82d8e2cdbadd72f317f86cf4fdf17af393e592cfcbcb;
// music[2225] = 256'h06d1adcf40c988d714f53dffb0ff0507ac07aef3e0de56dc5fde65e11eeb32f8;
// music[2226] = 256'hd7fb26f73dfcd8017501fe03be090d02e9e6c6dc6cdb54c8ffc076c1afbca0bd;
// music[2227] = 256'he9bf5dc294c2fcca62df6be3d1d3a0c2dcbe54cf99e168e369d82bccb1c706d2;
// music[2228] = 256'he7e2e7e283d168c3d4c631d925e439ddcecc26bdfebcbacb0cdbf0e0addf2ddf;
// music[2229] = 256'he3d3a0bd2cb244bc96d534e206def1dc1dddc5db19da09d83dcdbfb78eaeb6ad;
// music[2230] = 256'h3caac2aa0ba9c5a39aa2eea86dae17aa28a27f9dce9ee69ed89c1d9a2295b29f;
// music[2231] = 256'ha1b387bac6bb34bc58b66cac48af32c58cd375c95db788b1e4b4beb058a72fad;
// music[2232] = 256'h5ac09fc85ac6a3c822cda2c2aba1b78a7399ecafebad9ba561a9c7aca5abe0ab;
// music[2233] = 256'h10ad51ab18a970adcaae81aa04aa9ead3ab464b411ad86a897a53aa838b3acb6;
// music[2234] = 256'h20a5e290e68c388a9c876a989cb4aebf56aca68ecd84729556b15fbce1a6da8b;
// music[2235] = 256'h14870c91a19576942ba624be96bd3bb45bae8bae37b5b9b87cb800b373b372ba;
// music[2236] = 256'h9bba69bcdfbdd7bee4c0f0bdd4b9cabaa6bd1aab9f9972af5eca96d55bd02bbd;
// music[2237] = 256'h2fb7debc22bf40ba7ab579b88cbb94c1dcc482c328d088e41deb8bddeac59abc;
// music[2238] = 256'head291e764dafbcf11d39ecbe2c9c6d2b8d92addc7d8b2d0bcced2d7bbe216e1;
// music[2239] = 256'ha2db5ad64dcad6c338c409c23ec102c0bdbd98bf2bcf34ebbef642f0c6ef65f2;
// music[2240] = 256'hfdf14df96c024bf12bd942e0c4ed60ebd0e58ce28ae001e3fcf6170eab0e2609;
// music[2241] = 256'he80d3515bd16dd11c90f4512ba15c619131b771d6e1bf002dceb75f5160ab313;
// music[2242] = 256'h4517e61a8a1d11169701c6f2c907f12d1436dd30b63677352f27341611142328;
// music[2243] = 256'hc03ffe482b464c44703dda29ff199a1a182cb13e0f41be421c49bb3da728d921;
// music[2244] = 256'he3244e2dfa3ac538e320500d5d0b500fee0faf17932c3c39da2d9a1b7517a51c;
// music[2245] = 256'h4f1d951da929293d8e459c37eb205f1a861b78108b0a0a1aaf356443f22f9317;
// music[2246] = 256'h7914351a8f1ad01821269a37823bc73d7d4213462e4699469346da346c223427;
// music[2247] = 256'he1396a49ce43c42db0205a238e260a25a430394a6456cd438b2a0026ad28da22;
// music[2248] = 256'h711f1f3668602373656101433835603fb549a84bda55cb65c862cd4f32446a49;
// music[2249] = 256'h3c5e126e156d2c658b6226633e548d494a4a45370a22681f6025cc2d293b7e50;
// music[2250] = 256'h1155af3f4d29b5218b287c2f2d306838464c4053573d802632282d33892ed026;
// music[2251] = 256'hbc306741684b7c47fe38f62db52606226223a228f628bc2bb73fbc52d84cac34;
// music[2252] = 256'hc8240c2e26419f4bfd50f856f455a748043400253f22a1215724d835904f7e5b;
// music[2253] = 256'haf4a3c2f0a249a2779268f246a3349487b4d3d393f1ec417b91bc22107303647;
// music[2254] = 256'h6c5c65602c5d055cbf53e54144354f383139ae33352fd42baf2a8b3009490b5f;
// music[2255] = 256'h665a7d44b22e7031663e003e8e32ff1862088f0dc90fc60d3c1cc235883a9126;
// music[2256] = 256'hb00fef036005c40bfc14d3240434112d9412e1028b090720ff2e9f242a0c30f9;
// music[2257] = 256'hbb01a01e0e31ef2f522783250321b6104d07fd073205caffc6fa1afbf9021d07;
// music[2258] = 256'h1a0629023e08a31f1a285b1b390aedfb6df808f4e0f5cb07001b95214510fbfa;
// music[2259] = 256'h98f297ed0feb11ebf0ecb5eceeeee0ee42eca8f8ed0140fd05ff11105b22ae1c;
// music[2260] = 256'hbd099bfb10fe3511971a6019ce1b811ede16610d4b0e6e0325efdce785f328fa;
// music[2261] = 256'h25e513df3ff1e9f0fade24cc37c5c9c7fec8e1cbbdda9aee39f430ef7ceb39f4;
// music[2262] = 256'h72fe2bfbdcf709eb88e352e8a9db05d44ad141c451bd54ba91be6ec3e7cc05e5;
// music[2263] = 256'h2eec0be043de92e5bbde69c65eb75fc1ecd743e491d832c2d0b9b7bafcb447b3;
// music[2264] = 256'h08c7b2e3eee61ed100b816aa66b70fcee2d8fed95dd3f0cea8cf9cd58ed2fbbb;
// music[2265] = 256'h5daa0bac23bd0bc912cbacd7efe20de1d4d227c4b2c6bacebcd02fca83c1b2c3;
// music[2266] = 256'hb7c6d2bd99aea4a91cae9eb6ddc7dedae1deeccce0ba90b03aa1cf98dd95ed92;
// music[2267] = 256'h7c93e999b5a8a4abbfa31fa4b4a5809fc78e54846b8bad91ac8cc88b8b9f1db3;
// music[2268] = 256'h27a93391c48941918494e990478b2c8841874f8d0ba257ad4baa34ae78ab7f9b;
// music[2269] = 256'h128b8f83e6882089f387b39d2bb8d9bef4b936b333a9d198fa8d9c9531a6e5b5;
// music[2270] = 256'h68b6f1a06790cc9281a0a3ad04a8eb945189798a228d8d8a6494f1acfab32aad;
// music[2271] = 256'h8fbbc9cf20ca6ab5faa651ab6bbf08cb28c17fafb9aa36bcecd55ddec3cd89b3;
// music[2272] = 256'h19acfcbfcfd733dc77c44bae71af42aaa7a124a393a1baa112a2c2a259a444a1;
// music[2273] = 256'h8ba403a9e7b129c968d82dce3bb122a2a4b3e1ceaedfa1d5d3b919af7cb2edb5;
// music[2274] = 256'h4abdc0c4a0c72bc471be66be12c0f5c0d3c409c96acbcbca3ac880ca29cc11d0;
// music[2275] = 256'hffe4e2f29aec2fed79f3bdf683f6b0f113f1bdf359feb101adeb36dd17dd3cdc;
// music[2276] = 256'h57e0f2e337e635e7f9e989eeffe931f0a707e60f75095910e0244d2e21288225;
// music[2277] = 256'hcb270d2adf30a0333930aa29e322ac2a0a3276243b12ba117e254e330b358e37;
// music[2278] = 256'hfe38f9380f2bae186016f00cfffd710587150817fe170923cb28cf236c1ecb1d;
// music[2279] = 256'hba15ee041001ab122328342781248f2e8d2d962b0f2ce528b3284f291a30bf33;
// music[2280] = 256'hfe345e2ebd18b80f1d139d16bc14a413b326a637863aa03957395c352b24db18;
// music[2281] = 256'h6c1b941bc0161e1d2b345941d9401142d446c63cff20fa173e212f27b0273b2d;
// music[2282] = 256'hac399537b0368b39bf35f3393a3cc34a3c5c255c6a5e4a51743b8e3b4c4dda60;
// music[2283] = 256'hef5ece4b5b39623c4253535f105af9490342c351fd68d172a0690c557939e735;
// music[2284] = 256'h5751165c904abe33e32bf439a44f68571d46e42e4f25ff37e7575662015e1559;
// music[2285] = 256'h6e567551d94ff657034a673506355137ec3a063967318631a836df3a9139b839;
// music[2286] = 256'h3e3a013a3a3a37329e2d4734d33c6640fe3bf8396e3cae39b635003689360b36;
// music[2287] = 256'h4b326e33e43d0040114163406234813f6d59e65d23584a55885171419c2c582f;
// music[2288] = 256'h1849c5569d53265e77685865c068976c5c70e17053647b5a8a56e454ae572157;
// music[2289] = 256'h4251a74a59480a4d705346531c4bb145874d9d4cd233e522e4211720c724382b;
// music[2290] = 256'h5c22f2114f10b81c8828fa2673137c058f0631099d094b0b701cf428001ecf15;
// music[2291] = 256'hc015dd1bb324052667267e208a19dd1a951cf91e171fda1ef12150201018f912;
// music[2292] = 256'h7917ba1a401cb61e541f8425fa22191c901bcc06d0f046f28df5f8f5a5f6bcf8;
// music[2293] = 256'hb5f805f75c05f818911ab20b87f91df9cf0a1812c00c9d107115f2125d1bd329;
// music[2294] = 256'h0b2c812adc2d7b2d1f292126b6230422ef1d2e1b541eed205723da216519ae12;
// music[2295] = 256'h15148b1b0d1518023afe6a021503ca052e037eff45fd09f081ea68f18beb1de0;
// music[2296] = 256'h9fd848d7aade19eb8203bc0d31fd4bf4c3f653fd3403feff8dfc11fcbbfbb0f7;
// music[2297] = 256'h83f239f3d5faff01a9ff4cf96cf321f164f354f770fd0ff268dff8dd7ce05bdf;
// music[2298] = 256'h83daf4df8bf2cbf7c8ecdfd86dd3c6e6d2f5b8f670f3adf3a9efa9df6cd56fdf;
// music[2299] = 256'h49f354f78fedc0e80dedfbf385f16dee4bef03f65d09ee0f6d07f10262028009;
// music[2300] = 256'hc50f530c6006f5fe6aed6ad9dbda62ef3403560759f6c8e233ddcedcfdd71ad8;
// music[2301] = 256'habd650c567be1dd535ed40ea95d285c23ac322c382bc9ec149d5a4e19be2ace4;
// music[2302] = 256'h35e577e354e4e5e117de75db31daeade6bdf48de96e168e668eca7dc4cbe3eaf;
// music[2303] = 256'h34ab86b062b996c1fec49fc11bcdbadbeedb92db20dda5daf3cc96c13bc340c2;
// music[2304] = 256'hd3bd90c1add3d8e25cdad0c987c11ec754d527d985d7f8dcb5e05be12ce0e1d7;
// music[2305] = 256'hbcd536e02de6e0e112e2a6f399fd71ea5ade9dee6b01a50551014c01ea00acf0;
// music[2306] = 256'h2fdd29e1b0f75e08eb05a7f053db19dbd6ed75fed5fc29f01ce1f0d27dce92cb;
// music[2307] = 256'h88c663c7bbc3fec9c3e546f44af4e9f7b2f547efe1ea3ceae4ea0bebddec56e3;
// music[2308] = 256'h8ad258cf05d303cf61cdbadfb5f655f7c2e176cee0cf72d4bfd11fd091ceaacf;
// music[2309] = 256'h2cd079d3aadcccdfe2dc7bd407d896f311046ffc21f6c9f698ef89df69d833e6;
// music[2310] = 256'h5ffbb9fc8bf426fba004e505e30130f48cdcffcaffcb13da38ebc0eb62d940cb;
// music[2311] = 256'h72d1deeb3ef78aeb2bf1a4ffd904250a2c080200baf91bf77ffa5efe32044005;
// music[2312] = 256'ha1f352e2dae5d9f9fa0b2c0411ee27dd73cac9bf2bc6bbdaabf428fad8ed13e5;
// music[2313] = 256'he9e1bedb5dd0fbce87d06ec89ac36dc253c181c3c7d34bee59f160df46cd5ac8;
// music[2314] = 256'h2bdacbe63ce55fe58fe5a8e75de9e0eea7ef08d8e2bf4dbc59c38fc70cc6fec4;
// music[2315] = 256'hbdc128c7cadc3aea66e134ce7fc700d677ea18f0f6e0e2cba5c206cf9de306e9;
// music[2316] = 256'hace4e8e785effbe41cd116ca37c4fbc1e8c43dc4c1c305c667e5650e970ed800;
// music[2317] = 256'hd0fca7f7daeb87dd3de0c2edc6f766feca0151056df925de9dd3b4dce8e12de2;
// music[2318] = 256'hede3b2e315e34dd8d0c401c093c34ac3ebc1edcc50e7a8f078e08dc905bf56d0;
// music[2319] = 256'h4be3abe645eca1f620f9d6e78acee4c5bed138e61aeb99d87dc88dc640c7b6c5;
// music[2320] = 256'h5dc753d655e869e6f7d349c46acec2e9d4ee4de460e06edf11df16df43e86cf3;
// music[2321] = 256'h72f43ff16ddc34c085bdb0c665c82dc66ec45ac58ac930d79ce9adea77d6dbc3;
// music[2322] = 256'h92c177c51bc896cbcccc0dce00d437e4f6ffab062fedc2dd70e0c1e157e426e7;
// music[2323] = 256'hbee66ee322eace01700c8308d709b008b309ca0d490ca20157ea70e4bcf637fc;
// music[2324] = 256'h78f420f116f775fee6f3a9e1e8de3ce1a1d770d1c2e1b5f8acff6fff5c04f3fb;
// music[2325] = 256'h49e019d26ddca0e645e3b6e245f6be0a380ddf0c8e0a30fac7e489dc73eb4300;
// music[2326] = 256'h4c086f0be7107c1420041ae760ddf0df0be437ec5cfddd1bfc24bf0f6dfde2fc;
// music[2327] = 256'h87118b27de27891415006a03561bc02da229ee147f049c0a91237332402c5216;
// music[2328] = 256'hd205190fe71e5e2fc03a0631a528d92ad42cfd2c6c35d4481d518c4623337229;
// music[2329] = 256'h8733bb433e4f14487f3827300027a422df25312d682934163b14f41cac1df51b;
// music[2330] = 256'h8d173d19391da21a4f162f134117d61fb9246e21d41a201a881a381cb71cc718;
// music[2331] = 256'h5323893b5d47de394823ba1de51e2a1df525d22ea52e192884214d212c20c92d;
// music[2332] = 256'hb748974d6542c43761319e32a6357b364036ff39ed39c532ca3111393e438043;
// music[2333] = 256'h3a3c0f35522d2330db36df3b743ba836493d1038af227317fb1614198d18f92e;
// music[2334] = 256'h4d4f46536e54a35c565d915731533155eb488832cf2c423d344e224d594b4c50;
// music[2335] = 256'h4153f455a458dc5aae5b9f58534528319232e736ea3543355f361939c938d738;
// music[2336] = 256'h2637ed371636da27322034289e353038262b731eb61c412b313cca3c5a36173a;
// music[2337] = 256'h433fa332a4233420b01d24188816f726ba3a603d8d3bcd39b1356c33e8359a3c;
// music[2338] = 256'he43fda3cba365432a835093eca41cb4086390b2f0236033c3f2edb2665209b14;
// music[2339] = 256'h69163e1edd23a325fa24a0250d236c2b543ed83bc02ea731b437be3fb3514d5a;
// music[2340] = 256'hca4fd23dac34503dd1461647de4c445428542750db486747ce4bf74fc751294e;
// music[2341] = 256'h6852cf4d1937a931c02e4d1a9b0c1615d82c7739de363531df2d932e902f1934;
// music[2342] = 256'h102a4714231387148910b413e2162a1a8e15080a7b046e040d0d53147916b323;
// music[2343] = 256'ha82bff226c226628532bcb2ec62dc1279520af211e28a6286029e91b60012afa;
// music[2344] = 256'h4502ca07630a5d12642147260b1f6c1b041dff19e20e31083c12ef1b321c5220;
// music[2345] = 256'h5225812843291f29ee281d1d381f8830e5296518f414ee212631533560376634;
// music[2346] = 256'he62c4428cd2a42300b2dfa27371d1c09b3ff330d4824482c882077ff93e258eb;
// music[2347] = 256'hc2022b10fc06abef37e368e0b0e424ec95fb9c0931021bfad8f9edfe53033504;
// music[2348] = 256'h26065ff707e92cea31e601e186e5d9fa9e0c3a0c6709b00af40f5710e00f2106;
// music[2349] = 256'h2ae87bdd41e597e804ed7bebd4e3e8da40d8dcdf45e3f0e48ce5afe168ee0607;
// music[2350] = 256'h5f0b4bfdfce8f2e0fef45805710099fc3c05ae0d6cff48e75ddf48ea14fd7002;
// music[2351] = 256'h3cf0b5df78ee9808f5119211c710d4159612f600eff43ffac30ce9112a0b5f0a;
// music[2352] = 256'h3709390a15076b031a0496030a0890ff11e92bd6a2cb58cce4cbb4cd90ce5eca;
// music[2353] = 256'h80d738ea08ee11e173cf3fcc96ce14cdd8cb1ec94cc5ffc3e2c0d7b99ebf1bd3;
// music[2354] = 256'ha8dd81d134bafbaf9bb403b8bdb32dba71d262dcd8d566d25bce6bcabccae5ce;
// music[2355] = 256'hbbc8a2b0b8a558b637cdb8d4afcb61ca1fcd6ebfc3b04eacefad4fb18abae9d1;
// music[2356] = 256'h77ddb3d40dd0cbd02ad348d252d0fdccc1bed2b539b8d3b7f0afe3b6dbdcc3f1;
// music[2357] = 256'h54e4d8cf65bddcc4c5db38e1adde79e132e6acd97ac235be28c611c7abc433cf;
// music[2358] = 256'hf3e2e7e428d3c9c2d1b9ecbb8acb42cda2b4f19d13a26fc040d4ebcc56c80fcb;
// music[2359] = 256'hc2c643b887ac86b5bac611d160cb11b6e9a931a929a9c2ab42af03aeb4a540ab;
// music[2360] = 256'ha4c207cc40c019ae15a61fb13ac483cd00bfeea946a8f0b0f8b363ae98aabeae;
// music[2361] = 256'h94b07fb0fcb2fcb66cbb56b7a1b1a3c1fcda95da9ec907c517c8c8c776c663c6;
// music[2362] = 256'hb4c3b6bf42ce53ec7af807ef0ae628e3d3db2cd79be2c2ea41e9cfe939e6bddf;
// music[2363] = 256'h85d654d269d785d9d1e8cbf873f54cf69ff8a3f983fa2af7fdf72cf442f834f4;
// music[2364] = 256'hefca2aafa8b4d4bb9ebca2c0b1d205de49da08da3edcaad678c774bb6fbe29cd;
// music[2365] = 256'h11d9c4d496c546baf3bfb3cc65d28fd991e09edebdd762d834dd6ed1adbefbbf;
// music[2366] = 256'h77d2c1dcd8d8bcd5d4d7bbdcc8e105ea99eafbd040b6a8b7bccf7ae66be3dbcc;
// music[2367] = 256'hddbeeccbd8e6f2f4aae8f9cd6bc416caa0cb49ca38cc26d5c0da63dc4ed906d1;
// music[2368] = 256'hfbd771eaaef3b8efc1f41e062dfe14ed45ed8befbeec0eeabff92e0ea70ff00d;
// music[2369] = 256'ha2106912210500f5d6f5d3f049e9d5ee03f5fff840fac0eeb3da6ad861dec4d9;
// music[2370] = 256'he3e8a806a9121c16641905198015c4121e13b40aa3fa56f6000126112a18d309;
// music[2371] = 256'hf2f6b4f8930f8c26ef24a40c40f60ef6ac0df121f51ef30cbcf8faf939128c20;
// music[2372] = 256'hf021c5236524c122c91fad21a522631f3322eb1e8e0c9bfee207f51e1d2a242a;
// music[2373] = 256'ha82dce31db24c40d880a181379162a177111f60a480df5142917a41489111b10;
// music[2374] = 256'h421d472a2728ae27fa2ae02c5a2e882f2d2eca316d42604a3849004ec44f8e4d;
// music[2375] = 256'hcf4cce50a14cf6348525572c3d2c7e14510f902c1d3706256c0c43fb2e0a4723;
// music[2376] = 256'h0d27c424b9264e29252c482c8a2953269926382bcb2ceb29b22724279e28e027;
// music[2377] = 256'hec27b630c0326f20940bc20a4d1de12dd5304b313a320b24760a74024414d02b;
// music[2378] = 256'h0d37d428720c7804460f77135c0f610a66047d03e2199236fe39fa36b53aef3a;
// music[2379] = 256'h373c0d3cde365e313030e332e433a532772fa22e4436cd40ca405034c32a0025;
// music[2380] = 256'h791f11268d388a44bf398825dd1f1d24ce265923931b251741185725b63b2c43;
// music[2381] = 256'h323e154438428227c20d15053112262aea30e32e84325333ec307f2d482f9a37;
// music[2382] = 256'hb23c013cad34ee333a39042a5019ee1f8c306f40b03e3c2e2e257221601d1819;
// music[2383] = 256'h5c23c63ac23f9238b839453ce7325a1e58186b278836d1365b239a101a108e14;
// music[2384] = 256'he011db0c4719cb313e35f52be02abd2cb8306833bd33be346037c634b21ee70c;
// music[2385] = 256'h120e120f1a10540e660ec30d5b0c242a56481441452d1a21b025f5303a364e2f;
// music[2386] = 256'h581c6b158b157e1251139a1404151e13c51bee2ec33169213b0e560bd6118313;
// music[2387] = 256'h1617d0163e138f0fcd0841096007bff712eab9eeb4ffad08100737047a055a03;
// music[2388] = 256'h83f700f4bbf675f2c6eef7e95be718eb26efb4ee7ae7a5ebd1fa8e01b004750a;
// music[2389] = 256'h650c08f89fdc9cdc7de530e70ae534e03bdccddc1dedf7f86bf5dff9a101f2ff;
// music[2390] = 256'h05eb4cd7ecdafbdee3ddcee3d6f9a60d850403f2fbe3a8e843fc76029d02f002;
// music[2391] = 256'h5006b406d207121815124afa2df516007e161b1e9611ab03ebfcf10ca023cf28;
// music[2392] = 256'h2623851f1d1fbc15b5067f04a313e9227023080dbaed46ebfdfe380b94050af0;
// music[2393] = 256'h85e79fedffeec2ed6aec9ceb17e86beec803be0ee10d400e3010d0058af299ef;
// music[2394] = 256'h34f1b2ec75eb61eb01f0d9f320f4c5f2b7efd5fa710ab30a61ff18f596f5daf3;
// music[2395] = 256'h6aeefdebfbe6fcea93f39cf533f286e972e524e174e76e020c120e10870d9d11;
// music[2396] = 256'h141028fc87ef55f93d10221cd80c01f5b4e8bff6f30d7c155f16c013841a2626;
// music[2397] = 256'had27f521640be7f7d8f6adf6d1f452f6d2063415b6117f0fd00f5f10bb10060e;
// music[2398] = 256'hb20cf80dbd12b111c701e4eab8e4dcf320fc8bf155dca1d052d5a2db58e022de;
// music[2399] = 256'h16d856d5abd466d6b1d260db74f131f91bfabdfdabffcaf204db24d9ceea94fa;
// music[2400] = 256'h64f818e6c8d862d8a7e7d9f5d6f6aff5c3f31af73dfb21fde1f617dd77d1c8d9;
// music[2401] = 256'h82db6ddb37dcdfdba3d677db28f1f0f628f377f762fc9effd1fde7fabfefaedd;
// music[2402] = 256'ha2dd28ee2f025f0b7eff48eb6fdebbdb86d9ebda36ebd6f9abfa79f9a0f3eced;
// music[2403] = 256'h93fd2e0e170e22106d147411e9003bef1ff426066d13ad12ad0d720db3038ef8;
// music[2404] = 256'hbcf0dcea17f23ff85bf269ef7af6cef16ade15da1ddf73e1f4e087da1dd674d6;
// music[2405] = 256'h02e535f82dfa64f98cfa5cf9cef7c2f751f787e625d43bd956edfdfeeafbcce7;
// music[2406] = 256'h75d9c0d8acda58d782db38ec29f7f0edfddaf0d358da4fe0afdf26e486f3f2fa;
// music[2407] = 256'hc5f1f2e3d1df70ecd6f904f959f738fd7aff71f66ee7dee40cf20bfcd5fceff9;
// music[2408] = 256'ha4fcb8ff61f5bbedf6edf7ee6df5fff383f0cbf68efebc101c1fe51136fc1ef5;
// music[2409] = 256'hb3fb82fc1af756fd9f09cc0f810709f88ff320f33cf47ef94df26be065d81ae3;
// music[2410] = 256'habf77100b5f2c8e042dce3dd01dd76df90eefffe1afc97ebcddd22e325fa4705;
// music[2411] = 256'hbafd03f706fdfefe23eb4ed98dd6afd6f0d7cbe102fb1d09fcf7eae011d927de;
// music[2412] = 256'h10dfecdaa7e4f6f650002bffdefcaef8aaebb6df68e28ee8c0e194db10e779fc;
// music[2413] = 256'h4504a4f2c8e21ee0c0e0f0ec73fbb1ff3cfb4bf55fff27113013c70277f4fdf7;
// music[2414] = 256'h8a08461f1c2473132f0d170ea80a6f08800ef61f4b251b18980c6f0902130422;
// music[2415] = 256'h6d274c1efc0a57033a0da819d721ab1462f410e7cfee6cf02ef1e0fd1c0a250d;
// music[2416] = 256'h7c0eac11d50c6cfa20efd4f1b3f019eef1ed1ced7aeb5cea73ef67f048f41706;
// music[2417] = 256'h290bfbfd80ed3ae78ced9aee4cee1af064eeafecdbe898e934ee27f054ec3fe5;
// music[2418] = 256'h37e7ece717e6aff06d00a50850fff2f181f0acfb980ca804e5e659d5a7dc15f5;
// music[2419] = 256'h780011fdc3fb75fab8f9ddf8fcfcc1f88ce2e8d79fda14dc9ae363fae3127311;
// music[2420] = 256'h240a2f106e129c1246103c0b2b09d005b307600b6e0e38119e01e5eeb8ef46f1;
// music[2421] = 256'hdceca4ebe2eccbe817dc80d755d88fd2b0d1abcf71d463ebc3f660f276f012f5;
// music[2422] = 256'ha1f329e024d637e283f4defd4aee4dd704d037dd57f24ff844f737f6e9f23ef2;
// music[2423] = 256'hc2f160f54cf994fd3ffed9ea0ad55fd6dbe9a7f4b4ee96ecc3eb5eeaeaef31f6;
// music[2424] = 256'h9efa29fbd6f9c3f474e5bedb25e52cf7b7fff5f35bde00d982df86e0a9e0e2df;
// music[2425] = 256'h96df10dd9ed9fddb03d9cae4e8f8ccf90f05d8121a13cf145a18ba1f2f13f9f7;
// music[2426] = 256'hcaef19f255f625fb4608911523118b0b8410201d3b271229d91de1054afc73f4;
// music[2427] = 256'hcde80fec3dedf4eb23e9b6f0760b6711dd08ab07a7065f04140168076508fef6;
// music[2428] = 256'hefecdaf4690335099408c70a33082bfa55e88ee43eef06fdb501bef469e63ee7;
// music[2429] = 256'h8ff7cf03d0fd63fcce02c4fd67eac9d6cedb1bf5af040a038cfed30051ffccef;
// music[2430] = 256'h4ce2a2e833f644fe7d03bd080e0c94f9eeda25d890e442e8bfeac5f00bfd1804;
// music[2431] = 256'hb3f9faeb22e376e402f4d1fd0afe16ffa7fc06fcc6fa29fb240ac415bd12b806;
// music[2432] = 256'h0ffd61021a033cfcdbfd2e081517a91293012a00c4f9c9e486d95fe2eef52f00;
// music[2433] = 256'h48f8fceab2e71df0d7fd790109f42ce75ee591e945e98fe9f7fb080b3c093f0a;
// music[2434] = 256'h190c210b46094907eb0534f974ed4ff038f0a9ef10f984065a13ce0dd0f57bf0;
// music[2435] = 256'h0e01cf083c0871106f1f6226cb1a440afc08f90ad105b305df098a0ce40ac006;
// music[2436] = 256'h6606450a191ec933d42f4c1fbf0c1108b31a382ba63296322a3025291c14cf10;
// music[2437] = 256'h07253e384b476b42922d71258029de2bad28a4273a334640e038a02762218f26;
// music[2438] = 256'ha62aa125832923383440bb41a63685297d24db210c26a41f9d10970d7409dd03;
// music[2439] = 256'h12057108cd09ef0f3526b33a6237181e4206ec056b0e941118136a10bb0ae50c;
// music[2440] = 256'h391e992d892698112908680b8e04cafbf6042b17d71f8a127fffa8fdc70dc420;
// music[2441] = 256'h3b21dd17161a331fe714cdfff3fceb104f2218254f1fd61d7f1c2d0e3eff5dfe;
// music[2442] = 256'hf803d206c50c8c18821f421ed21b121ce61556041401ce15dd1fc618aa1d4430;
// music[2443] = 256'hdd3ba832cf1f3c1c54208a1b8416da135612bc14651d912e5633aa24161abf18;
// music[2444] = 256'h0e1bf50edefad2060f1d841d9111b9fe0dfe63162d2a8d271110b6fb9cfafc09;
// music[2445] = 256'hcb1c541cf20a3efc86fd420c7e15ec0eefff0bfb68ff60f98af075fb96142f20;
// music[2446] = 256'hab1b581cfb1fdb163c075303be057b0064ffaa10452b1336bb271019e618471b;
// music[2447] = 256'had1d03227d222c23cf22701e831ff81f3e206028f02909295f2c4d29f6256224;
// music[2448] = 256'hf92369264b24172906365a3ae53d673ffb38db3d544b914ed344ea35f532d33d;
// music[2449] = 256'h3a492b4bcf3c8d2b7627882c8e306632a93d034a5944a93d0f3fe033a5256224;
// music[2450] = 256'h51207c1acd1dae234b272526d1247423011f851c5718a419af152cfd65f47bfb;
// music[2451] = 256'h0efafbfae5f8def5caf929fc83fc87f720f487f675f4d0ef67eb95ea68f5bb05;
// music[2452] = 256'h8a0950fbafe916e74afa8e0cb50c160a370a1408d903d4fee9fe8e034807d905;
// music[2453] = 256'h63ff82f9e9f78afc49038cfe21eb97de50e71df7b1fb72f520f47cf4c6f13bf7;
// music[2454] = 256'h2efa8afce208890d200aa00b330a8cf962e89de79fe805e755e75ee96ae8a6e4;
// music[2455] = 256'hfef3d6043302f5025c07680ab008380548fe06e584ddeaeb13f1b7f6bbe8fbca;
// music[2456] = 256'hf0c358ccebd2d4cfebd333e505ed82f19af28fed9af03bf249f1b9f5aaf894f7;
// music[2457] = 256'h80eb84d94cdafbeaa2f44af2b5f075f54ff25ce3f8d76cdc67efd1fb58fad9fa;
// music[2458] = 256'h20fc8af7daf4fdf891fc8efbc3fd05fb0fe8e4d731deadf1a5f91eee5de00ce2;
// music[2459] = 256'h71f425020cfc6ff468f91d0084fc7cf507f3e1e52bd64cd7ead805e0edf40b06;
// music[2460] = 256'hd515f217d602d2f021ed62f2e7f368f567048c0ce20bc80f430f8b0ca80a590b;
// music[2461] = 256'hc609e6fac5f50dfb5be953cfb9cab9d30fdb49dea1d6acc7d5ce3ee77bf2aaf3;
// music[2462] = 256'h80ee6ae1f3d11ec27fbfe1cd30dffae4a9d70ac704c2c2c26dc0d2bf25cf31e2;
// music[2463] = 256'h9ce39dd3f5bd48ba3bcbdad8e3dbebdc3be1adde46ceb7c247cbebdcdbe38ae1;
// music[2464] = 256'h37e2b5e5c9e6c1e384e103d9c5c5cbbe41ca8edd5eea0ddf2fcdaec88ec970c6;
// music[2465] = 256'h87c19dc561c8efc433ce9bde9fe376d629cbefd638deadd547d6c5dc09df63e4;
// music[2466] = 256'hb6f2f3fe06f8b5e735e237e693e370d893dc92f27c001e021902abfe16f1a6dc;
// music[2467] = 256'h8cce4ecc68cc1ac7bec494c5ccc5ecd2b0e336e6d8e409e764e7d1dacbcbc6cc;
// music[2468] = 256'h3ecd41c93bd237e53cf2dcee64e91aed90ea25da2ecbc6c870c9eec869d1f8e2;
// music[2469] = 256'hddedeee640d819d17bda08ebffefcbe9fbdd40d89fe42ef49bf645f295f40ff5;
// music[2470] = 256'h96e594d448d800eecafd3bfaa6e664d511dcd2ef04fd1dfa88e679d635da23ee;
// music[2471] = 256'h9bfbb7f791e9c1d9d7e51809f8185d1041feb8f4f1f51ef261ed8df0f4f86ffe;
// music[2472] = 256'h3efec6fbcef67cf5b5f659f577fc5e0fdc19c00fca008ff10edeb3d95ae28ae5;
// music[2473] = 256'h31e7cbe86beab3eb46ea6dea0ee741e210e21be374e7eceac5ea1be76ae216e4;
// music[2474] = 256'h02e77be94de601e92900dc0cb80bcb0ae806800a990d060d07087704940cdc03;
// music[2475] = 256'hf7f0deecdcec17eb67e9f0f9600fae0f4f0b4c0b490fb814b81424125d0f680f;
// music[2476] = 256'ha91277183418c9133312910f1e0f5b0d6b108a171416661330044bf0c7ea52f5;
// music[2477] = 256'hb616552c5f2b4f2f7e31352e882abc282c20140f2b0a4916f92a5632e4249014;
// music[2478] = 256'hae0e8c1a61255c25492ec43c353cc92be4201a1ebe19d818ee1c2a20fc207122;
// music[2479] = 256'hed21a821f723b2222d234e19c1053002d907a5095209ef1114217422861d001b;
// music[2480] = 256'hde1a0e174d0c9f0b150b3303e601d302450636099f0a670df00c27151d1f601d;
// music[2481] = 256'hbb20ab267926be27a229432bc1299923661f3e1f0924ec27a328682b6725d811;
// music[2482] = 256'hd7053a108722d727ac1bd2087f0579141d26992b891ad607e30c4b221b34e736;
// music[2483] = 256'hca328b307d30b230813283313f238b14ee151329ea38802fc3265b24091fd920;
// music[2484] = 256'hb020e0239721f91212112112b611e8090bf1b8e88df2e4f7a5f958f487e912e4;
// music[2485] = 256'hc1e785ef40f35af1f2eeebf0f7f69ef6b9f33500220be3055f02d906af072efd;
// music[2486] = 256'ha5f5e2f674f612f260edd8fb290e0a0de90bc709f0054b08290a200beb080d0b;
// music[2487] = 256'ha60a53fdd3f10bf49f03d51008175e19c1136e10560ea60c5c0d330c710c4b0a;
// music[2488] = 256'hc60634097d08a5fc01f638ff9f0b27189615d004a7020410c920951f950d4506;
// music[2489] = 256'hf60cf41e6427432199204c21fb1e0c1c661de818d50792ff5d037304d0f25cea;
// music[2490] = 256'hf200cc09eb06270a4b07e704a900fcfd65fdb6fd5806f60333f619f212f58bf1;
// music[2491] = 256'h2aeadce83cece4f044f12def1ef0f7f28ef846fa5bfd8aff0a019a136a207119;
// music[2492] = 256'ha9152c1a071a070a62fe0304f0116e1f521be80b5d023f0724160b1999152916;
// music[2493] = 256'h0819201ec521b9223f12e1f6b6f0350377172216570da30dea0bcb0ced0eac0d;
// music[2494] = 256'h850b4e048909d11f6d2c362654112ffc51fdd20f611df718360648fdf401d503;
// music[2495] = 256'h6c048d04a502c3fed4fa28fe2301cf09811be1182f04d1fd34027af764e61be3;
// music[2496] = 256'he9e472e43fe473ef2aff80ff86ffc0036b05fa044cfe4afe4a00ea016801d5ec;
// music[2497] = 256'h16dfcde096e0a1e35fe641e8bce382e5cefba9051d0009fd88fbaffcd3fdaafd;
// music[2498] = 256'he8f323e260dee8ebb9fc9b02c8f8c2e730e2ceee29fd8700cdf9d4ed1be828f4;
// music[2499] = 256'heb037804700115024a027a024e044702f0f10ae4a0e7c0f652041900d2076923;
// music[2500] = 256'h9e26e815be08570956183b2105229624ba2702212a11650c100db006cc05dc08;
// music[2501] = 256'hd306f905af0685085509c1fd6bf06aee44ecc7e710ec8ffb6008d706b4014906;
// music[2502] = 256'h7808daf8a7e8f9e5bce5f5e219e531f6c50549003ef2c3e7e2e744ed88ea1ded;
// music[2503] = 256'h59fc240562fd56efd9e6dded20fde400270216089c08280772048d038f030e00;
// music[2504] = 256'h3301700302051b05cbf412e0ece082f419053c02c8f017e629ecf0fa9e04fffc;
// music[2505] = 256'h3be8a8ddbae254e389ddb8db37e35cf3f2eb85d546dec0ec8aea0fe74ee3c7e4;
// music[2506] = 256'h64e4c4ea35fe6c03df033b089805dc0137fbb6f8f0fdf90222045ff202dd95de;
// music[2507] = 256'heddec8d0b5cb4bcf93cd26ca85c90ecafbca8ecb7acac9cf98e35cf2b7e9a7d5;
// music[2508] = 256'ha8c762c423c4e3c604d6bce850ee4ce95be844ea3de364d40ecd1cd920e44ade;
// music[2509] = 256'hb6e0dded62f16eef08eed3eb1ce4a1d52ad4b1e564f249f2a3ecf2e5eae5d0e6;
// music[2510] = 256'he3e3ece4d7e84bf0afeed4d977ca15c91fcb3ecec0d5fee7edf2fce866da12d9;
// music[2511] = 256'h1fe8a7f5f4f9e8f2fddef3dd1bf08af10bef2e00b613041a7219201c341fba16;
// music[2512] = 256'h0e0ebd11ac1136093c08181c92303e2e442cb42e9b2d9430f726901177fc72ef;
// music[2513] = 256'h79f9dc0cb9166a0ceef4f2ed5bf5b3f891f7d6f5f0f6bcf893f803f59defccf7;
// music[2514] = 256'h5d0e5517fe0b94fcebf4f7fb9a07790cf707cdfa7bf3aafa8008540ca100cbf2;
// music[2515] = 256'ha0f259007508dd0704078e078e0555f382e60debadecb4ecd4ecd2eec0ed93ef;
// music[2516] = 256'h03018f077f077e0b6c0abe0a3b0ac50b52034cf179effdf038eef8e8dee1a8dd;
// music[2517] = 256'h6ee1daf6b505b700bcf782ee02ee56f514fcd2fd5efbdaf681f4a201fb0d8608;
// music[2518] = 256'h00fcf0f3dafaa608b10edd0b580ec11204fe90e250d8f3dd92f0f8f868f47cf4;
// music[2519] = 256'h37f729f1f1df12d8e4e611fca60039fb5bf83bf1b3edd2f2aefa8501bdfd9ef7;
// music[2520] = 256'hc2f52af896007703340219fec6f0f8e95eeba7e526e0c2e39ee74be585e6c9f6;
// music[2521] = 256'h530427fe84f1adec48f137f4c8f2e0f7b0054516c714dd0480ff4eff64fb87fa;
// music[2522] = 256'hb608311b051ea71ea81f8e1c7a1c07207a237820e11e101ff921ae3093318b20;
// music[2523] = 256'h6616541c112fac3a41390838243c10377920de15e11eb823b7214324842fc535;
// music[2524] = 256'h572cc6225427f225021189017207481bb626e11b400bf202e10b401cd2220028;
// music[2525] = 256'hdf2b3d2aa8267824f425db225c20c81e0b15da0dfb0ce4095c04540ac91f7c2d;
// music[2526] = 256'h3128db166408430d131ff529e0236e14630d8e102f0f1a0c44151f26ea30a522;
// music[2527] = 256'h9205b7fdb901c3ff86fe7cff9c009101a90f941f7f1baa1752195a191c189315;
// music[2528] = 256'h1d180f0fc9003d033b0b8a171a165303b605d211bf0f9a0d5210e31302155511;
// music[2529] = 256'h270d8a0ce214782765302a22380e170970110913430ebf16fe23e62830264f1d;
// music[2530] = 256'h3916aa0b99f898f4fd04ba12ce15f31149139a188b0cadfd51fb44f8aef397f1;
// music[2531] = 256'h96f7affc3f006a0fa412610b9110b017681a7c18e315f30bc5f929f65ef934f7;
// music[2532] = 256'h8efa5308d71aa11e950ba0f49df28c02aa10b7127f05d9f928fb3efe83fb27f6;
// music[2533] = 256'h83ff0210aa106702b0f077f00f049014f4165011700ea70786f846f045f97808;
// music[2534] = 256'h180de909a806480d34170e0b4dfd220572148d20ca1baf0c6e077104d2fe4afd;
// music[2535] = 256'h5cff2a02a904ae074705b2fe8e071b1a331d4a1159fb4fe6abe2b2e623ead9ed;
// music[2536] = 256'hc9ea66e9c7f7ae07a3023defabe23ee5fde874e48be837f91c06130215f1c2e8;
// music[2537] = 256'h6ee965ea24ec72ebf2e663e3e9f0a005db088a052903320332056604d403c3f7;
// music[2538] = 256'h5fe8d6e6bae676e4b4e7aaf87d0807063f055908ea01eaf29de561e864eda5e9;
// music[2539] = 256'h85ec58f9700168f68ee662e4dce700e7a7e0f2e346f59afce9faa2fbe9f7c6f3;
// music[2540] = 256'h7feed5e8c7f4a0073f0ed20f0b102e0b5bfcd4eb31ee3bfe260b2b0a5cf9bcec;
// music[2541] = 256'hd5f098ff7b0c3a0846f901edc7e35ce89ef779f299ddafd7bcddb6dfb0db07dd;
// music[2542] = 256'he6eaaff536f111e4c1dd94e74ff66bf979eb17da97d58dd922daf3d9e0e725fa;
// music[2543] = 256'he3fab7ef50e4e5e647f221f132ed24eb17e80cea17ec5deff6ef99ed0deea2ed;
// music[2544] = 256'h2af13bf143edd0f161f419f87f059b0dbf0243ed5ee62fed54f1f1f1cbefd0ed;
// music[2545] = 256'h02ee85eeb9ed5cedddf8630def1191ffcdeaedde66e3adf66f015e0aaa175d16;
// music[2546] = 256'hb516851da11b7b1a76195018ef18e5149513d014e018cd1eac1cdd1c2016fc00;
// music[2547] = 256'h65fa6df6b9e479de82eb66fe50057cff41fd5cffa80010021305c2fd7deb35e3;
// music[2548] = 256'hd9e25fe2a4e40ef0e702a6031ef4f6e699e755fcaa0196f41ef6d6f6c6f1f6f2;
// music[2549] = 256'hc6f400f7ccf546f43ff764f811fa8af3b8df18d86de496f4f9fc95f629e826de;
// music[2550] = 256'hfce2e7f3a6f8d1f110f4d1faccf4a6e189d736df1cede2f500eb5dd9a8d68ad8;
// music[2551] = 256'hc5d732d681d6ddd793d76de60eff1b0a0a0be9075007c809dc0a1e0d730b4e0c;
// music[2552] = 256'ha70955f6cce997e928ea84eceeee26f0c2edb8ecf4e96ee510edc2f21eef20e9;
// music[2553] = 256'h1de030dee1de4dda52d6c1d667db32def7e2e4ea96eda5efbdf47bf6dceb42db;
// music[2554] = 256'h5fda36ebc2f96efb52f9caf96bf811f8d7f959f23ce0bdd5c3df88f204faf1f4;
// music[2555] = 256'h0af1d0f4a6f6c8f53efa09f474e381e0e2e6b7ebf2ec34f4be03820542fe41fe;
// music[2556] = 256'heeff1ef754e6a6e5fbf4a8056c093bfac0ef50f365f9dff62ff36afe550a2812;
// music[2557] = 256'ha71441160d1ecd1332055309000b1106cc097f1bb92693244f250526e91b0508;
// music[2558] = 256'hc5fe940aec1bed220c166c0370fdd808c716300dd4f587e60ce2b9e2e2e2b9e6;
// music[2559] = 256'hf5e9bde760ea23f9a606a7002aed81de12e238f3250042fea5ee2be419e9f2f6;
// music[2560] = 256'h0e02aefd6af15de8d1ea24f98f035c00c5f1e8e91ce9bce4c7e64de83de915ee;
// music[2561] = 256'h37eea9edb6eb15ec17ec61e906f85a0c8412610e5a091305d8f3dfe4ade803ed;
// music[2562] = 256'h94ef3cf05aea6de74ee964ebd4e9b1e5fbe25fe1d5e6c7eeb7edd8f156fd0afc;
// music[2563] = 256'heaf9e5fe18f996fcca13eb1e7b1fae1fe01bde1b741e1b2102218b23c12add1d;
// music[2564] = 256'h28078f00640c7521b91b9efda0ece5edcf0024137413a811cf0e9509b311551c;
// music[2565] = 256'h471d531f43218e218f228821a1234b24f82129219324e22b7223a60bcdfe6908;
// music[2566] = 256'h6f1c3f26892bd630692fc529d12627273e199d0a1d0e280fc50e1b0ce5043606;
// music[2567] = 256'he80bc3132815671454245431df2e5b2ab72548237f265d29402ae42785242825;
// music[2568] = 256'h85261f2e8434a330612c3c1c6b092705e20786152a1d2521e433b13b503b3c43;
// music[2569] = 256'h7242e731f31ca6177d28343b9b40373f603ec63c8538c736d2355e2ac620b920;
// music[2570] = 256'hd31ecd1dee1ef5247825b5191c19b91ede1c2e181511c60dad0e2411a60b50fa;
// music[2571] = 256'hfaf2c9ff6a13401cf60f2df94cf26002a715d11b630cf3f8adf504f7bdf5f7f8;
// music[2572] = 256'h7307af160d17ce1426185617d10c5b039502af017cfbbafa5b0cd41c141e0020;
// music[2573] = 256'hc91d95182a1439121819111abd17400f6cfb30f786fb52fbc9f8a6efb1eef0f5;
// music[2574] = 256'h9cf97601a1061b030b06cd1194213e2fd22ca91ecd0fb30be4173123191fb60d;
// music[2575] = 256'hdf03960dc61ed22aa522590ff005600cc81cff2417257e1cd00e390f18147516;
// music[2576] = 256'hf513ab05f2fa78028314f21dfe216626d82665269d2378266c2be92c7b2f1722;
// music[2577] = 256'h1313bb16d31c1d203f23d1265f28c7259622971d7419c319d61c141fcb23ab27;
// music[2578] = 256'h7d2696250d202222b8315535ab322837423aa1303c1ac90a590cb811c212ce1c;
// music[2579] = 256'h262c9228bc1b3517e61a26205f22be1f0e0ebef53fef92fff612291757152d13;
// music[2580] = 256'he418f6260d2761227020a0197518bb1b4c20ec212a1daf1c831a6c0ec4049706;
// music[2581] = 256'h5311e21a94167808ea00ce0829167f0ee3f612e7d2e1eaedcefd05fd4ef7eef8;
// music[2582] = 256'hc8fe55f676e204dac6d74dd303d2f5def6eed7eea1ec52ed8cebddea0ceab4ea;
// music[2583] = 256'h55e95deb69efc0ebe7ebdde811d9afd235d937db4cd726d4cdd25fd3f3d1dcd0;
// music[2584] = 256'h57d337d4e1d495d45ed2c3cc0ac757d240e14fe08bd62eccd7cc04d8d6e24de2;
// music[2585] = 256'h83d44dc95dc878d78fe7a1e473e1bde051def0e14de525ecf1f6a3f9e8f14be5;
// music[2586] = 256'heedd6de334f14df874f81dfb56fee6fcd90071146f1e7d170e17b314b513d019;
// music[2587] = 256'h0e13ec06dbfd59f0b6e91aeec3efc3ec00e9afe6c9e968ec9fef6af02ef0d4fd;
// music[2588] = 256'hb4066d04c7068d0898087f041f0365002af3f9ee1cf231f430f1e0f193039f0b;
// music[2589] = 256'h840ec41619147d0fff097308d50b630fe314b10bbff88ff150fe4f1142154d12;
// music[2590] = 256'hc20d580cfb0cb60c8710fe0b6308720aa8fe3aeed7e993f5aefee6fdb1fe63ff;
// music[2591] = 256'h35fbcfede8e320eb9afe3b0cb10354fb61fa5d014e17e822811e3b18c815940a;
// music[2592] = 256'h8efaa4008afe7fec68e5aae188dfdadd26e8c4fae4fe03fd97fb21f9b6ec08e3;
// music[2593] = 256'hc8e57ad72dc9c2cc48cfaccb4ec8cdd2cce0b5e09dd63ecfa9d15ed17cd00cd1;
// music[2594] = 256'h57d092d132d10dd0f4c940cffce5ceee1ceea6ed24ed87e753d677d34ce3aff3;
// music[2595] = 256'h2af8a5e70bd502d391e45bf541f4d0f164f4d3f517ebefd747d3e2dc01ee1df5;
// music[2596] = 256'h6fe80ddf46dbd3d5d7d0bed619ee2cf9a3ef64e7c6e3f6e5d1eaf3edc1e860d7;
// music[2597] = 256'hb8ce43d70eed230422fec1e944e615e75fe438e480e886f03ff5b5f556f0deea;
// music[2598] = 256'he6f49003a90534fc1ef108f0b5eea6e81aeca5ec38e016dd34ecc4f7ddf217e4;
// music[2599] = 256'h17d6a3da99ec22f56ef498f2bef691f516e726dea5daafd867da46ddbfdf1eda;
// music[2600] = 256'h16e002f569fe2b0009ff09f9b8f3e0f81903bbf7afe43fe067e25ce442e7b6f2;
// music[2601] = 256'hfafc8bfedeff80018a00e1f305e7a3e53ce323e1d9e17ae594e720e8c4f370fc;
// music[2602] = 256'h72f6a5e8a8daa6df2af38afca7fb49fb47f9f5f16ee663e2e2ed5cf9a5026e0d;
// music[2603] = 256'hb910af12fc0c78fec0fc1e099d155b12c4023bfc05034112d81bdc1272ffdbf1;
// music[2604] = 256'h21f82a0cba14a4102b0dc8047ff55ce95ee522e64ce5c9e6ede921e7b4e2f2e8;
// music[2605] = 256'he5fbc80584fb1fee4be96eea50e719e659f4ac07b50b6afaefe787e43fe75aeb;
// music[2606] = 256'hf2edc1eb85ece0f0dff01bef41ed97ebc1eb15ebcaefd5f48df803096c12340c;
// music[2607] = 256'h5f0170f6f3ffe312c216a30f57087f0a93052df4b5ed3bf36ef54cf366f9a606;
// music[2608] = 256'h9a0fc90770f537fcd41149130312fc1fce280f28043532422140cb3f2d415944;
// music[2609] = 256'hd4453d416e40d63e0940933b772c5b2df1340532df2af921281f1f23ce2fad44;
// music[2610] = 256'h854f4945942e9822092dbb420b4da03e162c8a1fbd124a1125153d1cdc2bce2b;
// music[2611] = 256'h741d3f13d812f120812aca28f2261424ac26b22dd9337334a62d0f2b9c27251e;
// music[2612] = 256'hb8187d1c5f26db27bf21b22044261d25b9153b0e7510500ed80c910a6a09190a;
// music[2613] = 256'h600ccf0ea30c4e14a51fc61f1d175a0909077403caed34e3efe919e8dbe0efeb;
// music[2614] = 256'h13fb7ffe020160fd60f7bbf678fa0afe26f1aee7f7ec41edb2e674e59e00571d;
// music[2615] = 256'hda14b001d7f9f50474162a1a851c281d3b1b2f1cdc1c081dc3105cfd43f9b101;
// music[2616] = 256'h6b07e0096b0f75148d1215066f000d04d2f4a0e0d2dc27e94cfefefacbeb49ec;
// music[2617] = 256'h01ea18e6e5e530e41fe56ee3dee1d6e399e46bea4ef4a1f8adfcf200dffb9af6;
// music[2618] = 256'h8ff903fd33fc09f7d1f7a3fa48ef40ea08f3e3f5bdfb5f021801a2fc5ced4ce7;
// music[2619] = 256'he5f486f71df10aefd4eefaf2d9f4b6eb00e014e00cea10f47ef7c7f3acf28bf1;
// music[2620] = 256'h14ee6ceb38e6d5e192db47df70f2d9f9e0047e1b9f19a50c370cc911c719c61c;
// music[2621] = 256'h2822e029772524225520081f872529240228952ab619ca1b582c00332e2f851b;
// music[2622] = 256'h8011740fe8066009a4111015ba0e700696071c0d2c16f91aaf17750de504ad09;
// music[2623] = 256'h5a09e60c861de627c02ff628a31ec928e927171d5b183113ab15091573127b11;
// music[2624] = 256'h5fffb5f9d90be515301df317bf011301790e0c1247124b0d040463010b075b0c;
// music[2625] = 256'h040dd00c33104018bb16470966026e03ec08630e750eb90f6c136419be19d019;
// music[2626] = 256'ha52394188710cc2e523d8338893df03e5c3f383cb93f9a44c43289330545e43f;
// music[2627] = 256'hde3ccf3d8037b039a6427846563f4637ce2dee1fa920ce25d125f82b612d062b;
// music[2628] = 256'hb324f5182c1cfd231f2359218420a92415269427ac2ff02d2e279f2b4431152d;
// music[2629] = 256'h7f2b322d1d260f26dd2d113377333e282a2026213b285b300a2e34321c35c32d;
// music[2630] = 256'he62e4c301e2b6e22ea242e32a02fb0285925381f0f21d1259e2465200b1e4a1a;
// music[2631] = 256'h3113ee0dd1159529322dc826c12c8133fc31e22b492ffe320632903ba73aef36;
// music[2632] = 256'h9944a448e04829522d4d863e92381d2c8a275f38d340214b62520b421f3a8739;
// music[2633] = 256'h5132c8264e1e8923b61fd717091f8e214d1b0515bb13ef16e01850154b0c8809;
// music[2634] = 256'h780ebe13cd1ae719ef061af8fefaf1fd32046f0bb405cf058f12c01458083202;
// music[2635] = 256'h11005a00dd0e4613340db107e1fb73febb00ebfd1d0890059402f9070bf81de7;
// music[2636] = 256'h9de6c3e780edd9f2abe81fe502ee4de980e4d0e01fcc22c3e2c440b64db3b1ba;
// music[2637] = 256'h00b076b815d032d065d3b5d978d0cdcea5d452ce22c847d076d06ecf62d6e0cb;
// music[2638] = 256'h7cc576cc27ced8ce87cab1d1d7d56ebd20af0fb518ba3eb4f2a509a540ae96b3;
// music[2639] = 256'h1fb629b4ebac4ba8b4a969ac7db2beb0b1aa3db6e8c0b8c213c598bcd8b392b6;
// music[2640] = 256'h77bcefbdeeb762b7fec07bc1c0b96fbaeac050c748c9edc3fcbe95b9e5b6b4c0;
// music[2641] = 256'h63cdf2d044d21cd507d0aacab5ccadcd56ce79cc81cfc6d605d469d341d0c1c8;
// music[2642] = 256'h45cd17cfb7cad0c5abc48eca04cc17d7c0e9f3ec77ebe8ea1be8c3e4a7e3c9e6;
// music[2643] = 256'h12e739ec3bf6cdf85af683ef85eeafef07e4bae015e9a0ef06f159e0d5d4badb;
// music[2644] = 256'h94d99ad77edb0edb5eda12d65ddc85e5b0d67bcc92d55bd9e8d61fdbd8e21dde;
// music[2645] = 256'h01d5bed4d8d50ddd24e31fddbadb97dfa1e1d8e64fe999e178d481d2c1da88dc;
// music[2646] = 256'hc0e4fbee17df7bd1fedb4fe131e0aee5efeb10f08ff059ebc3e4bce651ed65f2;
// music[2647] = 256'h5cf96ef3b6e5b1e9f2f124efbfeaceeaadf121f622ec32e74df5df021e0c120c;
// music[2648] = 256'h7c015b0006fe90ff820f2a10cb07f10114fd5f015b028105fa08b0fb2dfbd20e;
// music[2649] = 256'hef0a37ea70d88edf69e455e530e970e9a9e81cf006f499e9d5e24cdf19dbd3e1;
// music[2650] = 256'h57e7fce652e145d914de6fe655eb59ec56e820ecceefe0ee8bf133ee2be21fde;
// music[2651] = 256'h2ae882e9e2e0c4e7e3f493f5ccef55ef09f0e2ebfaea57e986e652e75feb7ef7;
// music[2652] = 256'hb9fc36f93dfcaaf850ed82eefafa82fe72fa26f4a4ed01f73ffe6dfe430bc116;
// music[2653] = 256'hbb24df268b1adc1f3f1da21de72e2127741e6622931de91bb71fe924a7259e29;
// music[2654] = 256'h33310b21b50f7910d2085203970763063a0344fd95fabbf99af168f69fff47fd;
// music[2655] = 256'ha1fc8bfd2508cf10680260f9e602bd0cb60f05172322f72288223420771ffe25;
// music[2656] = 256'h4d1ccc11d8104f0b520fe914fe0fa208890869120f15b4116e0982fd9b038e0d;
// music[2657] = 256'h440c520bd00e4814bc150f19721be7170f1cfa1d011c10225e240528f833ff31;
// music[2658] = 256'he31e5a1ecf3d50537c4cb145c244d540d63dd838a335f03cee42a044f642c139;
// music[2659] = 256'h97356b32173385422d463d417a3d182b56221f2b2a2b7328832cb02d602d1c30;
// music[2660] = 256'h402b56285731e132322d8a2a5f29a72bcc2bc12764236a211026362a24266223;
// music[2661] = 256'h4223c61cbf1e942dc030d028fd22952180251c26c3239326c523e320922b762d;
// music[2662] = 256'hb3298a2fd926171a481b401f2b22b51b321ee92a9426e32399213715f716a922;
// music[2663] = 256'h0e275521b9224b338e374d3066342a3e3040f93bd83a2d39853568324628f521;
// music[2664] = 256'h1c25512807314e32082b572d68243510600b0f12381ab81b4815dc0a6d04760a;
// music[2665] = 256'h320f62101012140ce20aff10dd14ef190f17090956032408aa0b640bcd0aa70d;
// music[2666] = 256'h2f0dbd09a30886055e0998028aeebdf93310f9111211f40f0e09a3f9d1ebc1ea;
// music[2667] = 256'h9bf22cfbbefdae02e101cefb07fef9f60bf284f31dedc0ef69f073f164fc7ff8;
// music[2668] = 256'hd5f6acf719e82eee2e06bb0738feaff9fffa4cffe3003601defe78fe01fa58ed;
// music[2669] = 256'hb7eb98ec76ebc0f4e2fb66f720e0f6c141b943bee7bdb9bea9c7f1c4d7bbccc2;
// music[2670] = 256'h1dc7bac4e0be48b6a8bd3fc35cc096c243babcb598bac0b1b3b22bc14ac3e3c6;
// music[2671] = 256'h9ec485b839bb90bf73bc84b970bcd4c297bdd2bf9fc256b89bbcfdc26fc478c8;
// music[2672] = 256'h6ac204bb2dba75c45bcc0fc578bd27b917bd27c7a5ca10c6e1bf04c385c510c5;
// music[2673] = 256'h61c631c5f0d003e932f6d6f3def00deafbe1eff051fb22f522f863f641f5acf5;
// music[2674] = 256'h75ec4debecee88f5cfffd1fa75e72edba7e497f262f3d1ec8be6e2e86ef0c7f0;
// music[2675] = 256'hf2ed44ef96f399f73af3e6ec7cf65901c802f10091f8fef82ffdfff2e6f6d808;
// music[2676] = 256'h6607a5ffcf006fffeb0176079f079c05a5fb53f912036fffbdfda305e006b106;
// music[2677] = 256'h7907cf03dcf761f39fff6a05aa035009920e8f0a3607da03bafef204f4004ffa;
// music[2678] = 256'hc70dbb18e21da62d782d1525ae1d881c4321521b2519db1dbb1ce31f33289428;
// music[2679] = 256'ha22013202f21900ca8f288f6d30298fc1502e00d1a03e5f6aef5b9fba1fb51f0;
// music[2680] = 256'hd8edfde82ce06be355e732eb01f30ff751ef47e2fce288e850e65ee823eeaae6;
// music[2681] = 256'h65e182ea26e6dae39def46e8c8e5bbef92e7f7e065e339e610ea18e67de7efee;
// music[2682] = 256'h3cecbaeae9ec4bea1be467dd50e137eae9e9ffe875e64ee032eac9fc1f02f503;
// music[2683] = 256'hc70409ff06014505db05200a0b092d092c0f310dd004cd00f206ee04e8fde603;
// music[2684] = 256'h3bf911e9a4ed1aee8feef9eefbe9bde9b3de10da5ae45ce05ddd6be3b4e67fee;
// music[2685] = 256'h9fee42e62ee95befa0ec46e4eedf77e51de7fde61eedd8e5c7db7de1e9e64ce7;
// music[2686] = 256'ha5e77df119fa54edc1e5dfe882ea19f0f0ee93efdeed0de404e91de9b9e247e5;
// music[2687] = 256'h55e17cdf1cdfbfddb8e432e514de97ddeeecda03fb12611437088e0987130a0d;
// music[2688] = 256'h0d119320722728326439d8309e265220f71d872517216b09e8f96af4fef206f5;
// music[2689] = 256'hd8f6c2faf3fd6100e5fe36ff9f0040f888f36bf9b003ee0177f8bf0224090a07;
// music[2690] = 256'h7b0c890ea611510dff058808950ef61564128c14481c3b1632199118070e8914;
// music[2691] = 256'h7b20e627e429382384229529502a8826e72564295f2ce929db2dc2378a396630;
// music[2692] = 256'h842833283520fa2beb4d7b4f78451944fa426b43cd3b89401d4f2a53f74cce41;
// music[2693] = 256'hf53db4374e3e05494047944be93b3a2ff136bd2984201222c823bc254b24402b;
// music[2694] = 256'hdc2f0432a131282a4a23831eb3252f24ff1ecc261124932390217c193d1f2f20;
// music[2695] = 256'hcd1c1224a22ec12e7c26fb2008164414271ca618a81b0e1f47173519871a8316;
// music[2696] = 256'h3e1a0c1b401d1525df24da287333cb2fe41f831c6925b520a720ce35f444c54a;
// music[2697] = 256'haa49d940053b353b503daf3e28426241be3df33a4134b2327d309b38a8465735;
// music[2698] = 256'h75255f2c1d2a7320c61b7921d0263a23e01f7a1cc315e910ae17581ff41d2624;
// music[2699] = 256'h3329671f9e14e6134d1d491fe9100e0e8e13e70d8f12de162a106415ea156e10;
// music[2700] = 256'hc10a2503fe0b690e75061d06450093ffbd0169f93ff44cf66bf70dfbb10464fd;
// music[2701] = 256'h64ed59eaace25edfa3df32dbe8ebfdfc62f9a2efaae307dfe5dcaed7ded828dd;
// music[2702] = 256'h50e35edf96d17ad321d863d325d82bda03c665b522b9b6b8c7b8f3be0eb71db7;
// music[2703] = 256'h24be09b903bc03bb2fb09cafedb40cbc49c04fbd51b9b1bad2ba14b709bb02bb;
// music[2704] = 256'h74b9f9bf6abe4ebcd3bdbdbad5b8cab897bc0ec0a7c061c1fdc479cf2fd43cd0;
// music[2705] = 256'hedcc39c4d3beecc382c50ec6ebc76fc608cc32d00dcf7bcc76c207ccd0e548ee;
// music[2706] = 256'hdaedd2e96eea8deed0e8e6e4d4e05edfc4eaa3ef46e9dde8f7ec93f013f8d8eb;
// music[2707] = 256'h3fd0f8c960cf9ed9eede12d549d563d693d31fda20dde9dbf4d93ddc50e1b9dc;
// music[2708] = 256'hafd7c0d5d3d4fedb61e0d5df17e722ea6ce618e30bda3add4ce231d9a4e1fdec;
// music[2709] = 256'he6eb05f0dfe46dd53ae0b0eb4ee743ea5deee4e631e76ee9cbe89bf074f118ec;
// music[2710] = 256'hd4e701e5eae7dde979f4f4031f03e903ee0c440bb3047f01b0fd96fbf3ff7b08;
// music[2711] = 256'h410ccd0b1207ed00850be812390109f757f768f0f2f068f7cff4acee27ebbdea;
// music[2712] = 256'h03eea4f0cdf466f5ceea6ceb1cf37bec6ee763ec5df7abffe6fc84f5c0e95de5;
// music[2713] = 256'h1febffec69f207f789f416f70cfc80fd91f631eb42e993e7d9e7def2a2f147ed;
// music[2714] = 256'h2df8e3fb06f70bf3c0f173f8b0fb02f901f541f033f8c809100e690857076b08;
// music[2715] = 256'h180cef0b26060f03d9fccaff9c09d1074d023e016f0b22046eeb04f19bf704ef;
// music[2716] = 256'h24ed96e9c3ea3dedcdf04cf369ecaeec5ff2b4f510f370ec92f0a2f660f31bec;
// music[2717] = 256'he4ec47edcceed1f93df60ff3b7f864f66cfaadf370ea24ec16ec3401a00e5f02;
// music[2718] = 256'hdc042c0ad405a704f709180f250dce0bcd0c2912ac14d40d980b8d05fefea211;
// music[2719] = 256'h6727a2225a1a02211b23901d731610129217d11773154218b0162c195d1d2d20;
// music[2720] = 256'h631b7c10d0133d08e9fbca10fd12620ea9209425432577249219b316251a6a1c;
// music[2721] = 256'h961eff1a2f1737188b10f5012201ac0c7411150bc8096c0ab005b8079e0eaa16;
// music[2722] = 256'h161b0a1b171e231d7e1fb91fba1b892263214c2246290220d221ce2c052f1336;
// music[2723] = 256'he938c4341632d72990242c30173acf39383e9f41b443b645313fdc38ed378739;
// music[2724] = 256'hb7396d3f1647f93eb13c0b3f2c2c5f220a270d22f224d32cab283a2a5d2bd126;
// music[2725] = 256'h4b2cc5279e1d7427dc31cd30a72a02255224e325d3253f26fe29ee281a275f27;
// music[2726] = 256'ha125882b6e290925332cd82665210923c71fb7238325c020ab25702eb0264720;
// music[2727] = 256'ha62a83277e212625fe218d25a129ef227b1f8b29133546345c3e5647a3409f3f;
// music[2728] = 256'h1a349a29b12ee62a332ad22d152ad927e02a3e294a18ef0f19159a11ac160b1e;
// music[2729] = 256'h3b170015560dde02b10e7217730f890a2a08eb07f80c0f129a0fc00574024c02;
// music[2730] = 256'h7fffac02d103c4007904ab0aa80bd505c9ffd8040e0a7003e204a60b7a078808;
// music[2731] = 256'h8606acfef407a80abfff3904ea0e420ed2069e0509087b0099f939fe46093614;
// music[2732] = 256'h41150d0f380dc91264160510580e25156a158c10ab092e063e08a604f5fe21f6;
// music[2733] = 256'h5aea96e8e6e44fde1fe2d3e4b8e1f5db04d787dc5be47ae554e28cd8d5d096d1;
// music[2734] = 256'hdbcb17c3fec4d9cc2fd3a7cfa3c8dcc348bc49c3d6cc07c7c1c70dc309b92fc0;
// music[2735] = 256'h7bc4c8c202c21fbf80c103c065bb7bbc77bd6fc0fbc514c6cfbed1b8eeb6e0b7;
// music[2736] = 256'hfdbb03bbafc25ad53ddb02df45e0cdd877db3ade8bdb32da34d707d889d6bbd7;
// music[2737] = 256'h1adfb3dba5de5ce6dcd26bc02bc7f6cc0dcc48c74bc2bac6b3c803c962c959c2;
// music[2738] = 256'h36c641d2b5d496d34ecfd3c6f9bfbdc11ecb69d1ddd03bce8ed1f0d26fcf8ad5;
// music[2739] = 256'h17da12d988d8e6cf39cf26d878dd51ed08fb97f63bf5bcfb45fde9f9b3fa87fe;
// music[2740] = 256'hfafc24fecb0233009cfdcafd8cf783f6050cb921181fb117bf174f173b14b312;
// music[2741] = 256'h541710189a149e1459147e16e3153f16b31b960efafb51fe23fcb9f1fff64afc;
// music[2742] = 256'hc1fbec008a03040656022cf60ef6d400d506050056ff6504edf944f915037f04;
// music[2743] = 256'h3f02a3fc93019006e8044902b1f9d4fe3102befc0707a70a8b03abfd5ef9aef9;
// music[2744] = 256'h67fba300f305ce09910959032f027d004efe14047e0b73086505e00e260d7d06;
// music[2745] = 256'h340c720b3d07b8062a0b2b0b27012905bd08f301f2036a05f80561fdaeee1cf3;
// music[2746] = 256'h09f38aeb02edd2e952ed9fed78e525ed02ec1ee496e981e80ee461e02fe4b1ec;
// music[2747] = 256'h22e627e46fe508e0afe43ee64be204e666e9f2e9c0eb12e729df03e529e894e2;
// music[2748] = 256'hb6eae4f0f6e920e4dae1bbe870f4adf4dfec51eaffeb8bee99ee2dee2ef460f1;
// music[2749] = 256'h0eecc9f80e03db06b30644fd00012a092c06f80431025103e90498fba2ffad0d;
// music[2750] = 256'h620f7e0baefb97e5ace4c8ea38e66de9aaf045ee2eecb5e692e1a8e9b8ed4de7;
// music[2751] = 256'ha1e561ece0f226f12ee928e314e637e9dee6e7e781edbbf427efd9e2c1e363e1;
// music[2752] = 256'h5cda01db24dc41db6bdda4e825ee68ed9bf2edf34ef30aeec9ee9902ce0552ff;
// music[2753] = 256'h1c0aee0bd90359086b0dde0cfb139c1e6d239e203d18f6139313ff12c50e010a;
// music[2754] = 256'hfb0cd10d700be7106415b2132114ed0f71040905a20a2b0b840e3e0b1d036b01;
// music[2755] = 256'h480ae8104d079e08e2145519601d831a2b18301ade16e917f01cb01f27202024;
// music[2756] = 256'h1d2c972b3927622aa92c00235c20a72b122a9924222eba35a434363471336033;
// music[2757] = 256'h9839a5390335b433be2fb631cb2ff628392f012dcc2be841fa4f824b5c488f48;
// music[2758] = 256'h7a49164cf54c4d4a3845f4435045433d2a40a64c2c47ed44cb412034a4322e2a;
// music[2759] = 256'h611e7725be294f234f1f04237a26142658255b21ac1fab1f251e221cae164019;
// music[2760] = 256'hea1c3a193c1eef1f9a19bd19cf168e15311fdd23db1e371b751a57188218ed18;
// music[2761] = 256'hd9179e1fe72b9531a43274320231bf2d492c012dbc2eee2e612c3f322534912b;
// music[2762] = 256'h7436f6451e443446a446a13e1441bd469c41763e8740b03be23d5c4a21471843;
// music[2763] = 256'h934902398220c720e623081d5a19501edf21811bcc18ab19151bb221e81af60f;
// music[2764] = 256'h9910f60f0b141c179910ea0c5f0612fe4d02710fc311de07fa041306e5065e09;
// music[2765] = 256'h5b0a460ded0cc70d6b0d3b03080098fe95fefb059f0114fb75fa7ef580f216f1;
// music[2766] = 256'h89ef86f342f5e2edcbf494017afa2cf920f4c5e03adfefdf14dcdfdce7dcefe0;
// music[2767] = 256'h80df7bda27d5a7d06bd8a0d832cdc7c77cc256bcb0b9d1b791b5e2b2eab129b5;
// music[2768] = 256'hb2b7a8b97abb91b78fb7e1b98ab213adb8b3c2bcb6b80cb653bbfcb760bc39c0;
// music[2769] = 256'hb0b659bd24c4f7bbb6bcd3bfb3bbe9b89cb6fab88abe9dbf79c6c6c75fbd00c2;
// music[2770] = 256'hdec41abecac252c4e4be1abd6fc14ec7dec406cc2adf07e84ae7c5e0dbdd49ea;
// music[2771] = 256'h47f0f0e613e4f6e72de9a3e6f0e4cce855eaebf0acf2f1de63d511d9a6d7d2d5;
// music[2772] = 256'ha2d0d3d1a2d54ad054cfcbd0e6cc0ecc76d4acda6dd8cadb20dfa0db1ddb9cd8;
// music[2773] = 256'h77d508d9bcdbd5dc34dec8dbe3df6fe8fce170d86ad951debce588e41adf4fe3;
// music[2774] = 256'hd4e4bee73bee2aeb7cea55edb4eb76eaa8ea40ec97e6e3e3f3eabee5bfec0007;
// music[2775] = 256'h2f08d70061044d033e07cf0a4a05bc043607bb0794056f05740be509b5068703;
// music[2776] = 256'ha3f2d9e65ae5d0e896ed5be75ae8afec39ec7df338ee01e8aeed1debe0eb82ee;
// music[2777] = 256'h84eaa7e7c0e45de700ee7fef9df1a0f403f17cef04f06aea6cec0bf07bedbdec;
// music[2778] = 256'h8ce99fea22ef46ee6feb4eeb82f202f272eed2f54ff881f566f4d7f67cf9aef1;
// music[2779] = 256'hc1ecc8eda5eb28f846111213a007f60c9111570edc0dcd0962040e04a9095d0e;
// music[2780] = 256'he00ee00b960bbb12f8075cf4abf6a9f650eebdef8cef4cea18eb72edcaeea0f1;
// music[2781] = 256'h59ec6ee9eeec6ce832e7cdeab4ec15e98de175e748ec94ecd2f1ebec8ce73eea;
// music[2782] = 256'h13ef70f30ff2afee6ce8b1e8b9f05fee04eb6df010f04ceaf7efe2fd2107b00e;
// music[2783] = 256'h4e0fe9054101f904fc050e06f5076e08ec1325202a219129952a89235224df1b;
// music[2784] = 256'h4f16ed1c9d215223aa1e901d5620481ed91aca0bf3fb16fefe0353083e0b940b;
// music[2785] = 256'h0c137c1161ff00fd5b0a9a0fdf10a915e11e3429c9292b23d720bd1df418dd19;
// music[2786] = 256'hed157a11bf147c0eb106740a6c0f2a131d142e10130bcf0ac50d900e8a15261b;
// music[2787] = 256'h5316db138415481aef1f3d20561e271cdc1fe6279a291228372d623e514a6b45;
// music[2788] = 256'h0546c74f9750de44cb3776361f3b4e3c943cf13e5341a0429d483c462231b522;
// music[2789] = 256'hc32305281f2ccc2bae26fb23f9262d270a27022b02273025f82894233f24ea2b;
// music[2790] = 256'h292c592cbc2b2e29eb2bb12c112aa729f727192b3d2d2923ed22a7281224ff26;
// music[2791] = 256'h162ceb279326e028e525f822d126b8220923e52f002ae524a82c30260e214920;
// music[2792] = 256'h0e1b492397359f3ed93ca53e8b42a23f833dc93b9733b62d2f318732d42fab2f;
// music[2793] = 256'he72b722c932f5528c21f1a19311643169e154317ba12e3108d12c00b720b340a;
// music[2794] = 256'h18078c0ee70d240df61347129d0fe10b0106db07c8083505f204d3062409eb0b;
// music[2795] = 256'h2e0d2d0c5708480462045f067209460d7d0c7c0923081b059f0132013f07a30e;
// music[2796] = 256'ha90aad065d08f404690b32113b0eea1b69201119e51be912731024189d17e51c;
// music[2797] = 256'he717a0106514d612f9163b181111070ca5017bfb68fa88f85df4a5ec06ee2cee;
// music[2798] = 256'hebe49fde27db4ee0c3e449dcb4da18df31dafdd240cf08d339d600d1c9cee5cc;
// music[2799] = 256'h1fcb73c994c225c7f0ca5ec514c7a0c121bc46c089bd98bd3cbf11bcefbc4bbb;
// music[2800] = 256'h05b8fcb9bdb9c2b930c02dc12cbc78bc32bc58b91bbaa8c107cfacd7b4d960da;
// music[2801] = 256'hdad947da17dc08dd6eda02d9b5df4ee22ddcc2d9e9d89bdc8bddfcca7bc218c7;
// music[2802] = 256'h02c16ac371c758c485c3c3bd70c223c5d8bae1c0adc68cc339c919cafbc6ccc9;
// music[2803] = 256'hb7cb33cb79cc56ce37cf4dcf7ecc45cc85d114d519d671d340ce4bcceccea2d3;
// music[2804] = 256'h4ad52cd557d53ed4ccd3bad577e236f569f9d9f4b0f3f7f2c4f16df2aef766fa;
// music[2805] = 256'hbcffb0108118fa17bd1aee160714f613ab135a17e815b0147a184c18e1198c1b;
// music[2806] = 256'h84164e1053069afa9bfad3fd82fce9ff360247fd29f9bafb12ff48fee1017301;
// music[2807] = 256'h66faacfcf60158044503c0ff63ff0dfd8ffe8a0343047d031202f5066908c202;
// music[2808] = 256'h5c04c6050706c202f4fca002ea040904b6081605dd010f0746094f080c099309;
// music[2809] = 256'h4707810540073f091f0957120121e61e6b18791be31b441b691b72142607db01;
// music[2810] = 256'h780760051a0077011f01520138fca0efbded8ff017ea20e631e714e2a0e001e6;
// music[2811] = 256'h16e469e4caea75ec3decf6e482dfb6e695e7fce7a2ede0e95be84bec91ea42e8;
// music[2812] = 256'h41e987ea5fea2ae9dde72eea5de979e699edaaed3ee985ec34e6cee2bee66be5;
// music[2813] = 256'h3fe654e6c0ea78efc4ebffe9dbea2cf15df1faec03ffe80c370734070b066103;
// music[2814] = 256'h8209220bc60a5a0b2805b307770e5106ac005a07390908f907e939e80ae529e8;
// music[2815] = 256'h92f2d0f008ee67e769e030e55be872ea88e9e7e37ee5b4e75fe816ecb3e9b2e5;
// music[2816] = 256'h3cec05f2cff17ef1dbe92fe362e48de072e1b7ee63ef45e584e8c9e811e18ee2;
// music[2817] = 256'hc1df66db3bde52e2d1e76fe5a9e9e4fbcefc0eef59eb06f554fcbcf9ac02f919;
// music[2818] = 256'hbf248b22d722fd224b20041a2c175620db1ed212cc0f1a0e250e050cce0a1113;
// music[2819] = 256'h4f0a52f840f853fcc8fe4a0234ff12fdbc02c60624096e0b6008bf07bb0c8e12;
// music[2820] = 256'hdd133f10bc135a17d116071bad1d6320ef202f1f8623bf21671cb31b611f9e26;
// music[2821] = 256'hc0223621c5286c254c246527b026462c022f442a9d28062bba2a9d28682a4c28;
// music[2822] = 256'hf3265431353632359a40634964461347c8456345994a0c499e4cf94f3f479444;
// music[2823] = 256'hd64550493e4cfc476544b337a42abf2c542c122a892bd1272425cf275d255c22;
// music[2824] = 256'h4a25cc225b1c5c1f632bfe2b6921d5226d220c21dc261d1f161fde266c21e720;
// music[2825] = 256'h1e204b204325771f271c2b1e051ee41d511b3a1ce51c4e17c015631a1f1eca1a;
// music[2826] = 256'h1b17ef1f8b2c72313f30c32e1b35a2355b322841174c1f4d7951b94a5444b945;
// music[2827] = 256'h8d470b4ae142d83b013b633d03454f42dd3e90397c24e721052cb123011de21e;
// music[2828] = 256'h16213120e91793142a18c71bd71ed41f07210d1c8f16c51baf208b22da20af1b;
// music[2829] = 256'hd715520bbe0a2611ac0eb30ca90bbb0c820f930a170bad14c2158d10ae0fe70b;
// music[2830] = 256'hda0787094c067407310c8807c2053f021afc05fee2fe3cfca2f758ff8810c50e;
// music[2831] = 256'h930af50ed90ba10c0c0c3701b6004900f6eb18df62e457e300e0bde28bdaf3c9;
// music[2832] = 256'h12c337be43bb63c281bd43b6a8bbe4b778b9cebe28b711b6a0b709ba11bc7bb6;
// music[2833] = 256'hcab77bb6d5b292b507b734ba6fb728b46bb89eb788b4a7b2a0b4f6b61cb6f2b7;
// music[2834] = 256'h87b83dbb7ebd0cba24bc3dc1a3bf92ba43bef2c12abb8eba63bf51c1bdc071c4;
// music[2835] = 256'ha6ca54c513ce1ce1c5e031e3a2e268dc17df96dfcae6a3e9c4e2f5e3a9e1bae3;
// music[2836] = 256'h12ea3debb9f177eaedd38ccb24d040d34fd6c1da8cd5dccc68d23fdcb8d84cd0;
// music[2837] = 256'hb6d2fbd87edb1cdbfdd87cd993d9d9da2cdb6bd9efe0c9e1d2dcb3e1cfdef6d9;
// music[2838] = 256'ha1dc9bdd6fde6cda95dacadfeedb55de10e6aee2b8df70e1dde04de04de2e2e5;
// music[2839] = 256'h36e5c9e13fe2d1e1a6e390e777e500f01903340274fefb01cdfc6efc8204fc03;
// music[2840] = 256'hdb00a301a2007d01fb0425044705c60971ffa3ec68e738e8a0e83ded8fef61ee;
// music[2841] = 256'h19efb3f061ee89ea35e94cea55efd3ef72ed77f38ef611f5d1f36eef3ff24ef8;
// music[2842] = 256'hd5f3bfeda4eed6ef67f0f6f40cf519f080f11ff7b5f545ef19f04bf041ec60f0;
// music[2843] = 256'h3ff2d5ef0ef013efa7f094ee23e967eaaeed43f26cf215ef75f869059609030d;
// music[2844] = 256'h2b0f0f0f9d0c0f06e607630cd608a609690ad305b7026b08b90e92fcbfebaaea;
// music[2845] = 256'h9be326e9d8f001edb4ec25e82aeab4ecf8e6e0e914ebceeb6cee75ea70eafaea;
// music[2846] = 256'hbde8dce9c1eca8eae8e83beef9ec97e8a9e9e3e81aea75ebe9e8c0e86befebf0;
// music[2847] = 256'h8beb42f153f0b1e79becf1eb37ec27f341ee9cebdbec8af2fc00ce06490a670a;
// music[2848] = 256'h41067f15fe20571b031f07236e232e2686257d26ca22d51fbe216f1fa5207c1f;
// music[2849] = 256'h3822d72687138801f6fdf5f984f7c2f33df7d8fff700f6019e05d107260ab10e;
// music[2850] = 256'h9b063bfe4609800e571467216422d022ce1f641b4e1d4b1bd01a00172e127d15;
// music[2851] = 256'h2115280fb80a440c3c0f9a0f6f0dee08e50b380f35117e15b80f370d71151e19;
// music[2852] = 256'heb17cb160a19f7195c1d052d1f3db9416f4146450b472b44a946134d0850a84e;
// music[2853] = 256'he9516451453fda35a73ce03ea83a112d6a2138231524b1241e29442add29c527;
// music[2854] = 256'hc625a2280228bd25272bfc2a7b26112ddd2d6826b2299d2b7d29442ebf2c8729;
// music[2855] = 256'h892f9c2e1929e32bb52c6e286b29fe2c8f2bfb29e92a7f28d5220c21d6244127;
// music[2856] = 256'h1d27c7252d223022fa23b9222423a026bf26ab2017243735553e393eaf400e42;
// music[2857] = 256'h4b3e233c473b2938213bd83b8237fc3bcd3baf37a838f82e851f0b179517921b;
// music[2858] = 256'haa17ca14081a8d1cb6182a1538148b12d713f9152813fd1178138c15a9170712;
// music[2859] = 256'h7b0b560e3911bd0f090ef90bde095f0abc101012220d670d670953078d0c960b;
// music[2860] = 256'hd80cb30b640a1011cb0c4508900a700854093c09c9076d042cff2f01dc03f70c;
// music[2861] = 256'h9319fa1631171b24252bee26431f971ac214ce0e70107913f01327109d0d3a16;
// music[2862] = 256'h2510c7f5ebeeedf9c7fb39f7a0f8b9f62cee28ef94f004eec9ee81edc8ee04ea;
// music[2863] = 256'hbfe44ae7c8e038df68e028da95daffd82cd747d748d460d468cf1cc9f0c754c8;
// music[2864] = 256'h0bc9bac765c96bc93cc355bf96be23c248c7e4c5d7c08ac0acc015bdd3bd67c2;
// music[2865] = 256'h0bc4e6c38bc383c3d6ca12d721d646d2c6d85addcde1a9e0e6d61fd9d8ddf8d6;
// music[2866] = 256'h05d642dc55d7c5d275dc03d7bbc07bbe46c49fc2e2c313bebbbcc2c57fc2d8c1;
// music[2867] = 256'h65c5bfbfdabeedbf4dc261c7b2c6c7c5e3c4bfc4e9c615ca6acc83cc0acf44ca;
// music[2868] = 256'h60c3cbc6f9c784c9eac970c604cc83d2b2d2d8d1b9d115d25fd307d35ed078d4;
// music[2869] = 256'h48d7f7d33bd78ad7fdd15bd7b0e903f37bf10201e40f2b0af208b20dac101113;
// music[2870] = 256'h8215be18cd13040e040ec00d5f10fc104510481020098901bafcebfa49fef0fc;
// music[2871] = 256'hb2f818f6a4f6dbff440243fcdcfcedfbf2fecc05cd0093026e06dafed602c503;
// music[2872] = 256'he2fab9fd96ffba02b305f7ff54037e0333fd28ff6100eb0066fe1afc1c002cff;
// music[2873] = 256'hf5fdccffa0ff8bfdf0fb4afe0101bc0133ffe6fc23fff0ffcbfbeaf9e70dbd1f;
// music[2874] = 256'hf716ba17741ece1d0e23bd22eb214c228d20a71e751a6420bd19c005fb051602;
// music[2875] = 256'h58f3a7efecec97e6dce306e513e778ebdcecc9ea15ee24f07aec10ea02eecdef;
// music[2876] = 256'h63e867e712eaefe8bbeb59f03df282ec63ea06ef62ecb1ec94ece8e82ceca3ed;
// music[2877] = 256'ha9ef95efe4ea9cec1cecb2e951ec07eee3ebeee7d5eb7af10ced01ea7cebc5eb;
// music[2878] = 256'h40edb0e8dfe987ff530aeb05a809ce0ac20b6a0bfd048a09fa0c8f087d062502;
// music[2879] = 256'hb6ff1700d405ce088ff7d8e981ed63eb64e343e488eae2e8e9e4a6e9d9e841e2;
// music[2880] = 256'h5ae449e6f4e754eabbe9e1ee5fed09e317e218e89bee33ed83e968ee91f1f5f0;
// music[2881] = 256'hbcf14ef2cfecbae84deddae9aee65ced25ee03ebc2e726e3b1e009e386e4a7e1;
// music[2882] = 256'h30e2dae47feb4aef49ed29f8edfe02fb33ffce04560d9218c71d61218526a72b;
// music[2883] = 256'h812b46289623f01f8622071f20183d1eef1abd02aaf691f92ff97ff926f9d7f8;
// music[2884] = 256'h76f865f942fe95fea101ee01e4fc7903ec04a10181044e06ea0be30e7b0e5611;
// music[2885] = 256'h0615781611128614d91a3c1c421d151a0c1b151d9d1aae1fd0228420fb232629;
// music[2886] = 256'h2a291628c5274026b82bef2e4c2a552b242ae52c5534f12c7a2f7842184a4d49;
// music[2887] = 256'h2d49a94d2a50ee4b774e074f894b594c2546df4256443d45b44fff490d34992d;
// music[2888] = 256'h402d862dd32e932e6631492d0b2aa02d202b42281428b429f62885251c2d802e;
// music[2889] = 256'hfa243d26ff2441213c250824b8234a279b2534243124b920841da6206722b11d;
// music[2890] = 256'h5a1e76201f1c6f1b711ba41646171f1b481af319391a6517dd160f190817c715;
// music[2891] = 256'h131f5d2fee3d86423e3ff142ac4982469942bd461d4a684720456a462f47b243;
// music[2892] = 256'h7441de43913bba285c1f411f8a211b26922830258121ea22b621ca1ca21e9823;
// music[2893] = 256'he0204e1cc41e08209b1e781d781a4c1c5d1bb0193725ef251d1c671ed91a5b11;
// music[2894] = 256'hf8118d13bc10c50dc910c013a8100f110b1133114114d40ef50a490d4b0ee40f;
// music[2895] = 256'h7e0cfc06da031503660301018f0d171d8715c10d8d0e33108c12b910290f5a07;
// music[2896] = 256'h2501a405d90157016f0328fcd9fcbbebbdcae8c5cac8c9c58dc3f1bde0c06cbd;
// music[2897] = 256'he3b462bcd6bdb7b7feb8d6b7cbb5c0b75bbaf8ba4eb9f5b86bbabbbadbb875b6;
// music[2898] = 256'h90b8b7bb82b6f8b2d6b58db365b5e7b904b693b6aeba49ba46bb39be89bfb3c0;
// music[2899] = 256'hd7c1c6bc68bc23c59dc3e1be0fc085c186c7c1c894c749d499df89df39dfa2e0;
// music[2900] = 256'h66e37be327e327ea7aeb30e606e45be234e4bde4d5e76bec27db7bcab6ce9dd0;
// music[2901] = 256'h3ecf42d1eed3f2d31dcefcccafcfe8cd22cfd2d15acf6bcffed308d64cd3e6d0;
// music[2902] = 256'h4bd3a1d349d116d44dd70dd76ad71edaa7daead8a7d826d872db8add06d9f4d8;
// music[2903] = 256'h88d9a6dbc6e0eaddd3dc15e081e0e9e2b7e4e0e5f5e773e6b6e37ae48be52de8;
// music[2904] = 256'h00f48aff5f0093fe8001db04dd0090fe6e0379035e03ee055604e0048007bc09;
// music[2905] = 256'h9907e0facff051ee56ec2dee9df08bf016efa9ebdce83ee8bceb39ee9eed87ef;
// music[2906] = 256'hbbed99ea1bee37f135efefed75f0a8ef7aed50eeeaed47f01df19bedfded31ee;
// music[2907] = 256'h3ceca8eaa8ebc2ed62ea18ea65eed4eba4e861e9c4e9dfed45f10dee45ee2bf1;
// music[2908] = 256'hf4eeb2ecceee31f140f4a800df098405ff043d05300340031a01b307750c5506;
// music[2909] = 256'hc606190800077d05ed031b0663fc58eef4ef9bf1b3eedeee24efddf2c0f2f9eb;
// music[2910] = 256'hefecd1ed30eb53ed62eca3eb81ed4eed55ef36eeafeadfebcaed50ec57ebdfee;
// music[2911] = 256'h89ed5ce95eedcaef70ee63eedeebaaea55ecb2ec14ed4bee74ee5eedf1eb89ea;
// music[2912] = 256'h56ec20f210f2f9ebcfeae9eaf0ebc5eeb8eb23f28907e8170d202b21051c8017;
// music[2913] = 256'hbd150a18601ddf225c254e25a226bd24cd200b2447201b0c3a001bff55fd1a03;
// music[2914] = 256'hf1042fffbbfd25fb58f708f347ef81f02cf57dfbd6fc41ffc505f6094e0b5f02;
// music[2915] = 256'hb5fffe0d031312140f1da81fc01e592267221c1e1c1bbb1a251bed15f20f830e;
// music[2916] = 256'h820c2a0e300e440cb70ebf0d0f106e124b107e1596169f153d178d13341f9b32;
// music[2917] = 256'h9c353137a539293a293f8a3d3b3da944954328430848e3473246bc466b4c6348;
// music[2918] = 256'h9e36892c46256820182393224b25ac264621b323282666224e24b92564225824;
// music[2919] = 256'h3526d9242a29a22ae125c1257b273d28c12af72a1c285b27c828ff27a227ca2a;
// music[2920] = 256'hfb2b6e2924272227a929fa29d527c7270d270929a62de72c952d642e6b2a7329;
// music[2921] = 256'h042bbd2c042c5b31d140cb42843de93e553d523f813f133b9d3d833da83a533b;
// music[2922] = 256'ha03c6c3cc3386e3a9c37d224d61c90228920b21ef71d3a1add1ca01c5e181819;
// music[2923] = 256'hf716741535153612bb132117f7164614c012e7106b0e930f1b0e990f4312170e;
// music[2924] = 256'h25102811a40d0510bf10d00f850e1c0c480aec08c0081309370ba909ec085e0c;
// music[2925] = 256'hc10cd60ebd0d6c0b290cf7073a05da040f0ef31c0420ca1d151bca1bb71ae715;
// music[2926] = 256'h9119d41cdf207e1f6e19051e8218db111916690a81fae6f7b7f934f87bf63dfa;
// music[2927] = 256'h1cfdfafaf6f7fcf5fef49df4faf18fefeaf1a7f023eeabec97e8baea15ecd5e8;
// music[2928] = 256'hcfe84de602e366e1f0dca0da55dd8edb03d938db48d895d636d4c0cc0bced8cf;
// music[2929] = 256'h0dce22ccbec853cb0aceedcdbccb6dca9dcb66c73dc5cac1aec039d1afdc03dd;
// music[2930] = 256'h0bdc89d68fd511d6d1d27ad5bfd835d432d0f4d3fcd7e1d684d6c5d6a5cd70c1;
// music[2931] = 256'hb7bd87bea4bf07bf9fbf5cc064bbe4ba9cbefdbe2abe40bcc5bc0fbe49be65c0;
// music[2932] = 256'hd9c214c5a1c33cc1eac2c0c763caf8c690c7e0c861c6cdc85fca77cc97ce30cc;
// music[2933] = 256'hf9cd0dcf95cdcccdc5cf51d3fdcf8dce4fd58cd5e5d426d991d942d985db06dc;
// music[2934] = 256'h1adb6edf08ee7af886f6c9fc6b0ad30d6c0ba2086309ae0cdb0caa0b360b620e;
// music[2935] = 256'h67118a145415d207c3fdbefd57f973f95cfd99fdf8fa97f5e7f3e1f5d0f8ccfa;
// music[2936] = 256'habf9adf70cf7dbf9a1f9daf7e1fb49fca3f956fb5cfb1af815f71afba9fd8afa;
// music[2937] = 256'h45fbfeff2cfea3fb9cfdecfe25011e01cbfe15007d00160215045e03a905d205;
// music[2938] = 256'h8906840a2d0631035a054602a6086c18ca1c621d981fde1cab1cd01e8720ff20;
// music[2939] = 256'h941bb518401a731ad019d2179e19e2193d0ea104e2051e03aff670eefded4ded;
// music[2940] = 256'h41efa1f0a6eb73ec9cee6ce9ace7c8e55de53bea77e9b3ea3deb4ee86becb0eb;
// music[2941] = 256'haaea9eee2bec96ea7ce920e8b5e903e92fe96be95fe894ea8fed41ea88e6a0e9;
// music[2942] = 256'h39e949e693e883ecb6ee1eef36f2c6f0c6ee49f0d7e941f14705a1088f051b02;
// music[2943] = 256'had006a03f5012e02cb01ecfefc010d057e0418041804de053f0305f4e9e9e4ec;
// music[2944] = 256'h0eed25efaef23cee1beb27eb11ebb5e91ae973edfbed16eb7aeb92e9f6e7fbe7;
// music[2945] = 256'h91e5dae687e9f2ea8af0e9ed43e3ade477e9d6e85befb1f528f284f03bf3ccf3;
// music[2946] = 256'h67f2feee21edf3ec8fe90ee92bf09cf55af389efa3eb5ce697e53ce765e53fe4;
// music[2947] = 256'hd5ee0f001006f9069d0c1a12400c34ff8b05c00fa310cd1b0c1f0b1ec724d122;
// music[2948] = 256'hdd22cc1ed50e4605cd0046fef1fb38fa46faa7f654f361f280f407f85df72ef7;
// music[2949] = 256'h7cf83ffa35fa82f7fbfb01033a028a01a3027e020207210a300af3109b13e111;
// music[2950] = 256'h9116e0156c142b1b771d771c241e4721da238e229a239b28952c452f802e942e;
// music[2951] = 256'hd92f722d7c2f44323b3011394248844b5d49cd4810485c4a664ccd4933456445;
// music[2952] = 256'hbd4a2b494446924a034c8b4cde451536b9335b368a31753198316a2e0d2fee2e;
// music[2953] = 256'hda2a6f28af29d22c102ccd2702282527bd25c9286427762760298925db24da25;
// music[2954] = 256'h0827512964273226b72453224c24c7234c1fc01eaf215224ea245521ba1ebb21;
// music[2955] = 256'h70231422682589281824ae23de25472273216b200a2825358a3237351538a532;
// music[2956] = 256'h6b408649af4358433044de4686463c440445c245de46543bbf2c5f2ac0270e27;
// music[2957] = 256'h702bc7291a23c820cf20c71f371f6a1d052229284a25f92356229a1e2b1e021d;
// music[2958] = 256'h911c0e1cb11a081a631847180e17c8138e18bb22b921d81c7e1b3313330e780f;
// music[2959] = 256'h8f0cb90b240e771143135f13d6133f143f154012d10ff80f960cde0a2b0e381c;
// music[2960] = 256'hc026f91f851b321aa916b814b8133e14260e590b130eed08df062c0456ff9600;
// music[2961] = 256'h5cf503e780e71ee54de47de78ad70ec6b8c783c9b2c3bcbeb6beb4bfe7bf42c0;
// music[2962] = 256'ha7bef2be95bd8fba39ba18b85fbafdb9c2b402b7dcb710b7e6b7a7b76cb85bb7;
// music[2963] = 256'hb3b94cbb3aba12bc8cbae6b912bc06bdcbbd13bdd2bdcfbee3bf97c012c142c1;
// music[2964] = 256'hb6be9ac185c123c22fd3b4d95bd670d955d4fbd2bad84cd80ad9add8bed6b6da;
// music[2965] = 256'h32df01de62db19e106e2f3cf50c50dcabcc997caeacc4fca77cb46cdd7cddcce;
// music[2966] = 256'hd8cc43cceccddccd74cd04d0bbd0b5cd7bcfc2d0a1ce95d267d5aed49cd81ed9;
// music[2967] = 256'he5d51cdb77dddcd796daf8dddfdae4dbc5dd5ede80df06e22fe57ee3b8e29de3;
// music[2968] = 256'h56e35be5cbe365e29ce3fde2f8e596e595e749f7a9fe42fa2cfb79ff82021d03;
// music[2969] = 256'hf001c7fed8fc04000901ff018a022eff8a036302d6f015e78ee983ec3bed1eec;
// music[2970] = 256'habeb40e997e735eb0ded00ea0be776e6a1e8abec45ed64eb1eebfde9b9ea95ea;
// music[2971] = 256'hede89eec81ecc1ea5bed70eb98e999e8c9ea1af0a9eb61ecf6f146ec70eea4f4;
// music[2972] = 256'hedf25bf603f759f3dbf4c9f4b5f550f8e2f780f723f6adf556f605fb7607530b;
// music[2973] = 256'h6e06390742097f09e308180a960bca08fd08bd09e8093f0c360a440caf09ebf5;
// music[2974] = 256'h73ebedee51f03df2eaf287f27ef3ebf25af3fbf11def20f281f3b9ef8df0fbf2;
// music[2975] = 256'h1ff257f2caf128ee60ea21eab8eda3ecebe816ecd0eec8edabeed9ee94ec15eb;
// music[2976] = 256'hb8ecf1ec07eb57ed9befa3f059f2a9f13ef122efa0ed7af19df258f051f05bf4;
// music[2977] = 256'h0cf662f3c5fbdd08170bf207ed04da09bd0daf089712d023ca228e172a13031b;
// music[2978] = 256'he91d951c1c26d8208b0d1f0cca0f6f0b2609e407240492fe1afc5f03c708d303;
// music[2979] = 256'h23029a0014f9c8f620f767fa17ff52fc1bfae0fa12ff2f08ef0d7a0bc2011503;
// music[2980] = 256'hd60eb7117c17b22034229121791f3822b22634214c1c9e1b8c17971682172f13;
// music[2981] = 256'h8e11fb12b812df120c123810a50f411a002ac3298528f62db52dff2eba2ebb2c;
// music[2982] = 256'hc0308032813167337d374d38d939f83e6d36f429392a35290a2c6e318d2cce2e;
// music[2983] = 256'h10315223be1b351f38203a20c6218122fb23552852281c257d267d251c226023;
// music[2984] = 256'hae25aa25b726a62a892ceb2b722aa529d02de02f7a2f1333d4330c32bb31a72f;
// music[2985] = 256'h252e452ffc2fba3082328031f9310034b62e1e2c732e0f2e9735fd3f87441e49;
// music[2986] = 256'h0f4918461b442542bc42d43faa3eab405d3cf13b8b3d2f3ddf3c7b2e3520d31c;
// music[2987] = 256'ha1185f1c1e1f6f1ab81df21eb91acc190a17b616421b49193314f31432159d15;
// music[2988] = 256'h3d170d13cb0fda0fe10f8a110111a50f970d1b0d2a10e00e880f550fa109ea0e;
// music[2989] = 256'he513e00e540f7d11d20fbd0d0a0cb20b530d3f0ee40a510ce010280f490e9c0b;
// music[2990] = 256'h2a0f971e28231c2332256c20ee20901f391aa61f5520c01bce1edb1ced15c515;
// music[2991] = 256'h071d4621cf139302b4fda9f956f7b3f816f7c3f819fb22fa6df929f781f5ebf4;
// music[2992] = 256'hd5f4ddf5b7f450f575f861f8fbf4edeec3ea17edcbed3aeba1ebb1e8f3e4c8e5;
// music[2993] = 256'h3be1d1dc9cdc1cdb3ddd00dd2bdb22db3dd470d228d50dd056ce8fcef4cbe4cd;
// music[2994] = 256'h8acfcecd49cd3acbc6c4a6c63dd663dee2db91dc2ddd17de65dd79d7a0d6d6d6;
// music[2995] = 256'ha6d435d797d836d568d3cfd909da38c826bef4bf7ec05dc222c046c03bc36bc1;
// music[2996] = 256'h07c3bdc1b6bff4c338c5e8c4bcc3c0c225c45fc34ec3c0c406c507c3b9c3aac7;
// music[2997] = 256'h40c5c9c241c315c3dcc6f9c61ec522c8a0cbc7d029d1d8cea1d26bd311d14ad1;
// music[2998] = 256'h0dd51ed93fd691d5e5d708d4b2d3d7d9a3daced363d90feffff649f1fef0e1f2;
// music[2999] = 256'h9ff292f239f546f3eef355037a0c690b590bc7078f08dd0794f833ef4df43bf5;
// music[3000] = 256'habf466f7a0f4cef4edf849fa6bfa10f6a8f5ccfa20fafaf6fdf7b1fb52facffa;
// music[3001] = 256'h89fecffbbbfb6cfbbaf99efde7fd1afe05fd37fb48ff2eff6cff9902d1ff49ff;
// music[3002] = 256'h3e03f102cb004d03a804c8035c04c602fc024b074c0677010c05f006f5ff2309;
// music[3003] = 256'h351b9d1e0c1e481fc61e811c991a2b1b461b121c5e1d451da01a2617e7169217;
// music[3004] = 256'he80fa4fd89f639fcd5fee401c300ea00300101fb15fea9f8abeb41ea93e7ace9;
// music[3005] = 256'h38eb72e68fe835e920e9d6ea03ec96ea79e5a9e70deb23e987e85de7a1e653e8;
// music[3006] = 256'hcfed52f196eeaded61ee64ed34ec55edc5f1d3f1c6eef5ef26f097edf7ecc4ed;
// music[3007] = 256'ha5ef7bef12eee4f127fbf405f10804072b0add096c079706cd0485073f08ee05;
// music[3008] = 256'h48058602ed0295057202e5f55ee64be3ffe669e4efe314e94bea51e9bee99de9;
// music[3009] = 256'h65eacfe865e58ee50ce91fec94e96de855ea53e9dee96de9fbe8f7e9e9e72de7;
// music[3010] = 256'h24e520e517ea7feb12e9bae3f4e3fcebdeedddeb93ee9ff3a9f345f157f194ef;
// music[3011] = 256'h12f0fff0ddea6ce85ded28efc7ec86ea5feac3f3d5ff13ff27fb9ffb07fe7001;
// music[3012] = 256'haa00fa026d0ac91163117002d30251135e14611485121408dc0979096404060a;
// music[3013] = 256'h6109f9031a041d001bfb54fab1fa5cf9c6f591f50ef708f501f508f746f549f5;
// music[3014] = 256'hfbf94ffb40f9d1f900fdf7004d0379038807190f6c106a0e5b10c8139f166815;
// music[3015] = 256'hc3146019bd1bc81e382237213321d023e328f827b125402c2629a428ff3cec49;
// music[3016] = 256'h924a124b3e49cd478f474749a449c548a74a3447c546454d22483c4367467e3a;
// music[3017] = 256'h532aa1294f2b072ce42fdd2f062e172fe82f912d5f2bd02da62ed92b722def2e;
// music[3018] = 256'h422bf92a492d292dec2f5e2f4b28ca29e02cf8278128022ce5298627ae28392b;
// music[3019] = 256'hc0293027c927592778261627d727b328a028ef263e25d5222421f821cf1ef81d;
// music[3020] = 256'h8923bb1f18211e33c33a8639473d383c003ad43bcc387735c5368c34b0350941;
// music[3021] = 256'hb948aa47fb480d49d037f224ac2456278928442a3127b527b828de26eb255021;
// music[3022] = 256'hca1ede2030200b1e111fb31f741fa1252828182252209e1d3e19091c1b1dc118;
// music[3023] = 256'h6d16de19f81ebb1c24184e18b917c91ce324cc209c1cdb1b94162a15e512930f;
// music[3024] = 256'h110fa80c0c0e170ff90e9311a20e57133724ce2ad829ff2c462a592313216e1e;
// music[3025] = 256'he81c3a1b00185d1869144c100010680d8e0870f7a7e8d9e8fae579e6b7e799e1;
// music[3026] = 256'hfbe282e3f9dc5adb23ddf7d670c963c2f2c09dc063c258c0dcbfebc171be8ebb;
// music[3027] = 256'ha7ba69b87dba0cbcccb727b7bcb96abae0bb8fbaffb7a6b804baf8baddb9b8ba;
// music[3028] = 256'h83bd18bc9cb9c9b7f0b9c5bcccb8c3b9bebccfba26bf5cc08ac227d5d5ddd1d7;
// music[3029] = 256'hd1d9c4dbd5d9d9d937db60de50dc08dac6db5ddaa8dae4dbb9dddada4ac9f8bf;
// music[3030] = 256'hd4c3d8c2c9c4fdc751c5f2c455c60fc696c8a5cc94ca2fc8dfc982c936cc0ed2;
// music[3031] = 256'h93d346d3fbd239d12ecf3bd040d369d428d3c5d284d732db9edaeed8edd5ddd6;
// music[3032] = 256'hb5da72dd7fde28db45dbccdf22e1dfdfb2e005e49ae22ce2e5e4ace180e1d2e2;
// music[3033] = 256'h0ae3fdec42f8bffd10ff51fd85fe6bffb4fbb8f9e0fc9efefefb26fa8bfaadfa;
// music[3034] = 256'h55fa1cfce2f758ea1de4cde319e07de02ce3b3e2e8e284e48ee45ee7c0ebace8;
// music[3035] = 256'h97e680eb7fed12ecc2ebefecc4ed4ced1eea04e867eb3becfbeb42ef53f04ef2;
// music[3036] = 256'h43f41bf362f067ed73efd5f04dee92f075f423f4fdf3c3f498f275f362f70af5;
// music[3037] = 256'h6cf210f3d7f367f6f7f50df508fe8d0a4e0ef70d940fc70d6e0b610dc90f140f;
// music[3038] = 256'hec0b84098c08e1081f064e04890a28034df1c3f0a5f11feb92ea94eabbeb7aee;
// music[3039] = 256'h88ed44ecd9eaacec14f0f1ecdbeca3f0e6ee20ee34eda5eaf9ebd2eb54ec29ed;
// music[3040] = 256'h03ea82ec93ef9bec90ec10eea7eeb6ed5feb47ed67ee64ed18ef4eeff6eea6ef;
// music[3041] = 256'h32f033f1f0f116f4c9f246ef43f1dff1c6f1e1f1c9f04afc9e0ad50adb09220e;
// music[3042] = 256'h6410b20ed40c540c48091b08ae0a26083305fc0d5d1e901f850ae4fcbeff0a02;
// music[3043] = 256'h08067f08ff063f0994095a08ac0612041204710051fc0cfe43037f054200a9fd;
// music[3044] = 256'h39fd47f91af6e9f406f715f8e9f89afc3f007e06770bff0c820563fd3e07fb0e;
// music[3045] = 256'h3a11ee19a41cbd1edb200520871fcc1ccd1c8918cb1257134910fe0e8c0de10c;
// music[3046] = 256'h70199123a723ea230525c926dc26bc252b26e42414252c285e2ae02d032f962f;
// music[3047] = 256'hb531ab27681cb11e6f22f9234c249223f424af277a296828fb2af22d402f7132;
// music[3048] = 256'hd128281da9204f23c3228223ca223d22aa223c25d0267d263928472c702e752c;
// music[3049] = 256'h8c2c542e892ed52e592e342e412d3e2d662fc02ed52e0130aa30fb31e52ed62c;
// music[3050] = 256'hcf2ee82d662d362cbb2c383a65441d40803f9c40b63e3e41133fbd393f3a053b;
// music[3051] = 256'hcf39ce387f38d036c836d23528297d1e0d1f4a207e211320c61c6c1bf619201b;
// music[3052] = 256'h151b1e19eb1a5a1b9c19b21a4b1c361c2f1d241c8317fc160a179314dc15ff15;
// music[3053] = 256'h92149216ee1778160c147a139b13c2125013d812f610dc1036117910e0101713;
// music[3054] = 256'h1a129910f30f280c530ca10cd50aa50dce0a3d0edd1f9925b1227623cd24a725;
// music[3055] = 256'h3721bb200d236c1da01cfe1d511b4d1c6b1ac51910191b0a49fedbfe6f02040a;
// music[3056] = 256'hf5096103e3007cf90cf449f45bf1aef0f1f091f0a2f2cef374f487f493f3b2f1;
// music[3057] = 256'hd2f0bbf1b4f04ff0b1ef16eeaef071f1e1ede3eb33eb93ea7ceaf3e9b7e6e2e2;
// music[3058] = 256'h02e319e377e0f4e04ae146dd7bdce0db94d767d521d34dd2d0d1f5cc14d254e0;
// music[3059] = 256'hdfe250df83e0e4dd99d816d7efd76fda4ad963d6e9d667d642d5aed486d6f7d3;
// music[3060] = 256'h27c4d5baa2bef9c094c0c0be6bbf96bffebb2ebdc4be79be47c020c0b4bfb3c0;
// music[3061] = 256'h31c0fbbf81c15dc17ebffabfb3c1f5c29ac223c15cc2d4c48ec6a0c608c5ffc4;
// music[3062] = 256'he0c5b4c646c747c81eca69c908c9dfca4fcddcd0f9d1abd1d4d0b8cfb3d213d3;
// music[3063] = 256'h39d2c1d427d4dddb46ebebefecf11af31bef41f02ef0bbee2af36ef3f1f185f2;
// music[3064] = 256'hecf305f76df3bbf4a5fc5cf72cf3c4f663f6ddf663f67df558f6e1f485f365f2;
// music[3065] = 256'h45f3cdf40bf589f853f972f794f805f7f4f4cff731faa5fa0dfccefb1afbe0fc;
// music[3066] = 256'ha3fd8afeeaff61ffe3ff39019d01d6006fffd3fef5fe9201b403bd02bf026904;
// music[3067] = 256'h6006830425016d0285028f01b7ff16fe150a7a1780189218b31556128715eb14;
// music[3068] = 256'hfa11a512bf1363133a12ad1426152513a01654108b00f0fd690083fe24ff10ff;
// music[3069] = 256'h0cfeddfd8ffc96fc1afc94fbeefdf2fd81fd290085fa47ed5fe903eba7e832e8;
// music[3070] = 256'h7de8bae88eea70e915ea5cedffedf8ed1aedddece1edeaed6fedecebd3ecd6ef;
// music[3071] = 256'heeefbaef4bf0c9ef2cf12af35af010eec6eea8eceded2aef31ee60faae065906;
// music[3072] = 256'h2f055e028500e702ac038a0270001601a7010b01890320025501390240f799eb;
// music[3073] = 256'h61ead4e909e9d8ea3beaeae77ce7efe6b0e6e7e64ee5c9e4a4e692e7b3e61ce7;
// music[3074] = 256'hd0e78ae6a5e640e797e7a9e9d7e9e3e723e742e9b6eb4aeb33eb8eeb37eb3dec;
// music[3075] = 256'h66eddeef1df119ebcfe709edfaeea0f02ff558f58af570f431f389f409f15cef;
// music[3076] = 256'h46edb5eacdf61c040d063402c5fd08fca7f8fdf73ffa37f86ff85ffbf8fec203;
// music[3077] = 256'h7705f3098b0ec2fec9eb1cf224fb72fc4103ba07600b7d0db10bde0bcc075a03;
// music[3078] = 256'h49008bfb89fb9ffaf2f6fcf3fdf2a1f443f315f286f341f498f545f61bf7abf9;
// music[3079] = 256'hfbfbc0fc8dfd0400ea00de00cb03c507650aba0e38126411a91323163317151d;
// music[3080] = 256'h6d1d271c4a2047211e234c239c279d38143f9c3bc43da63ece3f9b415c413a42;
// music[3081] = 256'h3943a545c246ed464c48cd45c9464747833bf23322344632a4333d331131c532;
// music[3082] = 256'h4e3231327331592f1630f52c912c3330dd2c542bb82d942eee2ee72c792c7f2d;
// music[3083] = 256'h492dee2dc72d812d162f0d3194307d2edf2d6c2cbe2a8c2b782c882ba22a6a2b;
// music[3084] = 256'h422cf12baa296a28ae2a312b56290628e3275e27752467291e37223b01373837;
// music[3085] = 256'he7368d3545369d34db324332c4315c318a30ac321133e5348f348f245320b92c;
// music[3086] = 256'h542cf7295b2a64272b28a329f52b6a2c2828ef25312426220821991fcf1e371f;
// music[3087] = 256'h3d217f22bc202a2036200f20e5237f2486212d237f21b71e0b1f661bb01a611d;
// music[3088] = 256'h461dd31c4c1c421ca919f719e822c6240a1f841c5b1788120d11090e380dcf0c;
// music[3089] = 256'h0f124d1fac21e81fe3239622f3205a210f214d20d71c7f1b481ae4186a186117;
// music[3090] = 256'hc619a611bdfebaf6edf57ff30ff125eefaea58e89ce6b3e348e111e0addd2edc;
// music[3091] = 256'hd1d9e0d467d242d4fcd273c90ec251c146c013c0ecc07bc04cc060bf23bf42c0;
// music[3092] = 256'h19c096bf14bfb0bf73c1f8c02ec09bc0a7c017c0a4bf93c06fc0b9bfbdc04cc0;
// music[3093] = 256'h9cbe0fbd70bde7bd49bca6c3d1cff6d13ed176d2d1d28dd3aad34cd45cd417d4;
// music[3094] = 256'h76d5c0d58dd698d766daeedef9d67fc8efc46fc5e5c499c5a8c53fc663c724c8;
// music[3095] = 256'h55c887c8dec81ac9f1c9a5c728c651caa9cbb4cab5cbc9cb5dcc5fcd67cef7cf;
// music[3096] = 256'hc4d073d1abd1e7d292d5e6d5f1d419d6d7d7e9d739d84dd907d9e8d89dd98cda;
// music[3097] = 256'hf1dbdedcfcddb3dec3dee7de4ddec3df63dfabddb8e871f575f5b5f526f7a5f6;
// music[3098] = 256'h47f80bf84af871f9acf91afb88fa8dfb41fd62fd310061f8a7e923e870e971e7;
// music[3099] = 256'h9ce870e809e89ae84be841e8d2e794e871e809e618e60be681e4a9e566e7c6e7;
// music[3100] = 256'h84e81ce9b5e9c8ea01eb67eb31ec02ec25ed41eff4ef6bf04df181f29cf287f1;
// music[3101] = 256'h9ff102f208f2a1f29df34bf458f4dbf433f5fdf4b9f3b7f112f27cef71ee3efb;
// music[3102] = 256'h6f05e2033c046204a00399048a03e5031b0404041c057a040007fd07eb061c09;
// music[3103] = 256'hc2ff95f25ef269f222f140f232f1d5f08cf016f012f051ef3fef23ee91edf1ee;
// music[3104] = 256'hdaee82ede7ecededabeeaaee53ef58ef10f0d4f040f08ef0cbf009f150f245f3;
// music[3105] = 256'h40f43ef527f59cf491f410f478f362f3e1f201f38bf382f455f556f4c4f415f4;
// music[3106] = 256'h49f1dcf1f9f041f40a03030bf708d409360abc096b0a9b09a7096a09fc08ae09;
// music[3107] = 256'h6e0ab50bc909cb09ba0938fd97f3cbf399f61501a1026cfabbfd0b01b400ef04;
// music[3108] = 256'haf058604aa040704b703a1021f00bffc06fa37f87efbd4022f01b0fc15fdcaf9;
// music[3109] = 256'hbff7bff8cdf78af9f8fd1602ef04ff070c0d2b13be11d705e3055511d414e11a;
// music[3110] = 256'hd221d1228925f025bc23f11f051b60179a183a24a52833230323d7203a1f9a1f;
// music[3111] = 256'h101ee31f981f2d209a234c240226e626332866254d19da13fe16d9171d19491b;
// music[3112] = 256'h281c941dec1e69204122e221bf2235259226fa28892ac22be52b0e2b7f2ed92a;
// music[3113] = 256'h6920b31f8322d0224624bf241d25d52532270c2bf02d262e2a2ecb2e2030bf30;
// music[3114] = 256'h9630a1306b30d6316432ad31ca322532ad32ff32892fc82e452d2e321c41d044;
// music[3115] = 256'h1b42f5430a4388429142f9415a42ba41f54329455f432443fd408441093eb12e;
// music[3116] = 256'h5328192aa1278c27d1261c25f424f023d622e21fc41ed71eda1d0c208720df1f;
// music[3117] = 256'h781fea1b351a151ae1190e1b741bde1b291cb51b671b521a4719961af91b681b;
// music[3118] = 256'h6a1b761bc01a3c1a2a192819ae1859178e179a16b5148713dd1343169d145610;
// music[3119] = 256'h860d230a0811831ff1201f1e1b20d51e1a1ffd1f791e161e5a1fa524f0251023;
// music[3120] = 256'hfd22f91fe11e97193409fc0307086206c7054b05eb0272013a00ac0412093604;
// music[3121] = 256'ha60084ff23fb7af9f6f79ef553f538f3d9f2b7f49af545f7d6f7b4f78bf808f8;
// music[3122] = 256'h4bf7b7f7aaf6eaf454f5f9f404f3c4f129f02feeb2ec12eb1ce9bae6a4e42fe3;
// music[3123] = 256'h05e17fdf7fdef4dac0d9c5d7d8d210dbe9e6b9e55de46fe4ebe1d4e0f1deacde;
// music[3124] = 256'ha7dfcfde50deb5dc2ddc0cdc3adae3da25d33ec310c09bc21ac144c11ec0d6bf;
// music[3125] = 256'hd0bf6dbceabafbba62bc44bd61bc68bde3bd96bdf4bd68be33be49bc2dbdc1bf;
// music[3126] = 256'hefbf9cc08ac122c2e0c3eac4d0c5c4c746c87cc9c5cc5acdb6cc31cdb5cc40cc;
// music[3127] = 256'hb3cc30cd59cef1cf1cd0c9d0afd083cdfecda7d09fd082d0f8cf3ed012d280d4;
// music[3128] = 256'h17d69ad62dd7efd6c2d8e9d915da33dcaddbd3dc1cdb5add88ef38f9def738f9;
// music[3129] = 256'hdafadffc05fbf701cc0d920bdc09150cde0b590d460de40c230e0d0f3b0fa20f;
// music[3130] = 256'h190f140fad0e850d1211ae09c5f7c8f49cf7edf6b0f904fc8df866f6d5ff9a06;
// music[3131] = 256'h06050805610472053d06fc05ec06ff05f806e505f60450063d047206420a7607;
// music[3132] = 256'h34029afeb3fe79ff2400dafff8fd81ff1b03bc01f6fff0035c05cb04cb064c04;
// music[3133] = 256'he7019f00a0fc41fccf000d071b07e6fd97f749f8a5f8ebf83efbd3fb8dfc5ffb;
// music[3134] = 256'hc0f989fed8ffd5fdf5fd24fb1bf97cf793f874fc45fdb2fee0fe0a003701a0ff;
// music[3135] = 256'h4803fc0444085815911e302359251d2351212f1e8c19ca1a88200621731f2221;
// music[3136] = 256'ha420d01f271ec71857137b0d3a08dd077a0cfc0fe21121128801dbeb37ecb6f3;
// music[3137] = 256'h1ef290ee7fedb2f0c5f554f7eaf26ceef0eb65e73aeb86f585fb34ffc8f841f0;
// music[3138] = 256'h80f00cef3cf2d5f945fd26fcd4edf6e1d2e581eb72f7dd03bc0039fcf4f73bee;
// music[3139] = 256'h34ee8ff1baea98e4b2e6a7e9b1e6f2e788f085f51df7b8f30ff04eef70ebf6f1;
// music[3140] = 256'h35fb44fba6021a09ef05400259fcc0fa3e012203f1fc79f972facff53bed00ed;
// music[3141] = 256'h38f3def3a9f030f45ef754ee96ec87f809fb8b03071395134f1929237928eb2c;
// music[3142] = 256'h0d25731fce20a1238c2a312bcb2e84344434d733d82f692f0e314f31743ac643;
// music[3143] = 256'h2445714496436438182b852ac5229b19982717358635c43764359f30a235a837;
// music[3144] = 256'hbe35f835eb36653c51381430a836003d1d3f614256415236e029f62afb308537;
// music[3145] = 256'h5e3c693bf33e743f3d37d52c7f2cea38083ca73bd43d3336c62ed22cf92f4433;
// music[3146] = 256'h9230ff30aa32302dcc27322eb1355e33e32fb32c6f2ce52d14291223d020b325;
// music[3147] = 256'h112b192a00291c24a219a1142213e20b37071b09f809430aa00337fefffc3af0;
// music[3148] = 256'h9ef2720b7f140311bd0d320327ff3b089c0490fa73ff8102bd01a00239fd3cf5;
// music[3149] = 256'hb7ec70ed63f052e901eb6df1fcf51bffe1ff52f7fae327ccfcc851cf46d1c9d9;
// music[3150] = 256'hbbdfddd8b7d07cd1c8d4d9cfadcbc3d1b8d510d217d045ce89ca6ccd35ce49c9;
// music[3151] = 256'h81cdf0cf25ce46d296ce6bcb3bd028d04bd0c9ccbac5f1c2c2c04fcc63da60d5;
// music[3152] = 256'h9dd4ffd6bfcfaecf90cfe7cd29d3e6d54ade34e384d693cfcbd54fdccbde5ce4;
// music[3153] = 256'h6eeaa6e5f0e36de0b6d395d744e215e3b9e726ec93e8e0e407e483e278e7b8f1;
// music[3154] = 256'hdaed52e191e2d1eadfed36f09ff07ef79909f20d3f09d20abb06ac054f0e4c11;
// music[3155] = 256'h170bcc07ed0d2110a70c6d0b620bfd0e3413931a9125f620db15c617b41b3021;
// music[3156] = 256'hbe179aef45e2fcf522f93efed8076f08de0c080dac099b05db01bd024d023807;
// music[3157] = 256'h420df709f2fcf5f65503b90689010102ec03ea064ffee9fc6f076f0baa15ac13;
// music[3158] = 256'hb904dc032e042805a409550de814d8190d186115d61303120d180523cb245124;
// music[3159] = 256'hf5254b273d285f28c029e724d21f2a287d30182b0a23bc24b02e0c398a396c35;
// music[3160] = 256'h5f335d2e5c31d637aa357a3147308239893e15388c3b6e3e94321529b838854a;
// music[3161] = 256'hd14111453c564b547152f950814aac4b6b48ae458e4fb754b551ca493a403244;
// music[3162] = 256'h0249cf480a4f994b5342c13daf3eb7465d42233b3b39de318b327d33a4345338;
// music[3163] = 256'hc62cd226d62bdd29a02a0b2c581c3c062b0541104e12d210d80b8301e1ff3e07;
// music[3164] = 256'h7dff95f2eff5e1f22aef79f53ded6ce354e4c1e770e71edd21de00e442d6e6ce;
// music[3165] = 256'h7fd305d0faced8d375d3a4ce79ca60cad4cae6cb97d2ddd2b2cdc0cfffce16cb;
// music[3166] = 256'h37c876c01fba18bb84c3d6c501bc70bdecc6a7c820cfe7d3d1cc62cd3bd3aacc;
// music[3167] = 256'h3fc4d2c1fbc2cdc49fc777db00eef0e55fde27e107e4fce339dcbddcf8e2a8e2;
// music[3168] = 256'h43e85aed00e9f8e39fe388e58fe6f7ec7def5ce6ace513ef70f108eef0e936df;
// music[3169] = 256'hccd41dd329cfb3cf75d71bd881ddeee5a5e02bd8ded5ead8e2dc51d810cd5fcb;
// music[3170] = 256'h59d868e375e3c7dee1db6fdad6d5ecd285d7cedb83dc7ee11fe2ecd732d5d7d6;
// music[3171] = 256'hb5d699dec4e3dfe43fe5b2dbded4c2dc5ce707e63de317ecdcf205ef71e730e7;
// music[3172] = 256'hdee9f9e3dbe5c8e72ed6e5ccabd7f7dd7ddec1e8e3f174f25af886fa7ef7c0fb;
// music[3173] = 256'h96fc83f869f53ef14eec16ed82f2d0ec16ecbdf92af660ef99fd040de1164e1e;
// music[3174] = 256'h571bc811ee13ea250c316e2a8d25b32b9132323ce043ef3e7c3c793f513f3341;
// music[3175] = 256'h7d45e74bd14bb048784e6e457434f736ed39643e004c034a1d414a43b942a741;
// music[3176] = 256'h8f47c54686466e4dea47183f70414e430844ea43bf411b42f142c3442f43723d;
// music[3177] = 256'h773bd638dd350d3a8e434349c343ed3a1737083a163f953b3f3b3841483f863d;
// music[3178] = 256'h763afb38e73f2e3a8732923490321e33b23136350e3e1f34102f4d32212a672d;
// music[3179] = 256'haa37fb36aa30362abc27eb27812a6528de207b181e0eb30eab0f03078a044400;
// music[3180] = 256'h66f899f034ef4500770d4f109611ac0b2a091606570026043f061804c502e2fc;
// music[3181] = 256'hcefae8f925f249f2bdf5a1f75a006ffd32f69af2a1e489e2c5df98ce1ecf60d8;
// music[3182] = 256'hdeda39d5f4cc5acdfdcb4dcffdcd79c147c5f8cc01cc18ca76c8baca7cc5b9bf;
// music[3183] = 256'h9cc3d3c451c197c1a7c7e6c737c761cab4c8c1c661ba48b27ec03bc598c60ed0;
// music[3184] = 256'h09ceeec92ec55fba40baa1c65ccd60c9c1c825ca36c7dfc8abc966c884ced6cc;
// music[3185] = 256'hcec68fcba9c9d5c3c5c878cfa5cf0cc6bdc222cc9bcb76c18bc3f4d00fd496d2;
// music[3186] = 256'h77d5bbd074d029cf64ca71d567dad9dbf6e02ada5be6c8f4ace548e5c3f128f3;
// music[3187] = 256'h70fcf9fc6af132f52ffc7efedefe26f91ef3e9eed4f7c904b20597079703d7fe;
// music[3188] = 256'h8a03fd036b0810057aee75e2e7e14bda92d693de49e23be4c3eaf9efe6f823f9;
// music[3189] = 256'h04efdfef8df202f2caf86bf8b8eb79ef9af250e5acece9ee7de4bef01ef4a7f4;
// music[3190] = 256'hccf83bedbfefa3fa90fdbefc8af7cbfcc003e404da087c092105f005900d1911;
// music[3191] = 256'h251128110f12a3165c173a135011ef1c0e2df0312237a9355f2e572ac71f5520;
// music[3192] = 256'hfe2adf2c213138387b393b380f3a48393e33b02eb531273a6c38a437833b2c30;
// music[3193] = 256'hec368f516f54f44e0f4fee4d1c4e29483b4c1e5a9259a4584c51c542404a554e;
// music[3194] = 256'h274b5b50af4a044ac052d755b250843e3b3ec44bf442a5372a379733c02ff333;
// music[3195] = 256'h06394832872c5431942fd529932e4d2c8c1f92201e29ba22ed10eb0b5316e419;
// music[3196] = 256'h921afa1e7a1abc125b14dd158e106910ab0978f53bf294fb7efca2f994f4eeef;
// music[3197] = 256'hceeae1eafbf3c4f186ec08eb24dcdbd8dde358e189e06de4bde457e009d35dd2;
// music[3198] = 256'h5bd9a3d955de45db2dd3bad017cd86cedad2aad2e4cc25ca33d176d54ad37acf;
// music[3199] = 256'h03d16ad264c893c6a4cea8d3d0d596d543dfb8e857e70be8c9ea55f0b4ec60e3;
// music[3200] = 256'h49e87cea9bea2dedbae7ffe6b2e649e949f082e87cebcef8e4f284eee7e95ae6;
// music[3201] = 256'h7bf460eeb9d829d3a5cd81ccd6cf67d228dd3fdda9d7ced6d8cb04c65bc97fc7;
// music[3202] = 256'heac637caa3d251d936d37dced7d269d900df7ddb63d553d3d3d1bed797d95ad4;
// music[3203] = 256'hf3d5e5d51bdb49e0b9d81edbdbdb06d317d739d696cfb1d620dd25e159ea22e9;
// music[3204] = 256'h41de34dc81e2fbeab4f09fe92ddcdbd679dc03e5f2dc39c657c341d49bdb6adc;
// music[3205] = 256'hd3e2cbecf1f346f3eeee0eecd4f09ef546f1e3f05df405ef90e1e4decdf18004;
// music[3206] = 256'h1f0a2e06ea04a80c230ea80d99102d13da14b310d2126417c115fb1cdf252f24;
// music[3207] = 256'hb11ffd2264287829a12c4e31f938dd3aac287a16931c5a2a1a25ac218e2b8e30;
// music[3208] = 256'h133198292920931f2c257e31f7355931582e212ff22d9c27662c463785389b34;
// music[3209] = 256'hba32a131652b60315c385b339a3520359037a736a127392ddb376e325c2d732e;
// music[3210] = 256'he0324731062ddb2ba930003087294a2f6d29a221822a2d29442a502cda237e1f;
// music[3211] = 256'hd81b6c1b86221e29e228702847281520fc1ed91ccd16bd1cf21ba717791a4217;
// music[3212] = 256'h07109d09cd09a10ab7055708ca154d20ce19de0fc810f40cec06b8043eff02ff;
// music[3213] = 256'hb60445082907f802d4fdd3f4a7f2c0f792fbfaffb8fa0df30aede1e762f17ce7;
// music[3214] = 256'h64ce05cfd5d428d9eed77bcd62ce54cce9c816ce8ecd6fcad0c9feca4dc9c3c0;
// music[3215] = 256'h08c0f9ca83cc05c255c4d3cfedccc0c19ec24ec881c6f6c5e8c530c9e2cd15c7;
// music[3216] = 256'hc6c57dc5cdc061c62cc336bdf8c2eac38cc5eecabfc7c6c241c6e2c54cc4bccd;
// music[3217] = 256'h4ecb00c44ccaa7c352bb39c39fc201c67fd789daeed635dbe9dc85dc23d81dd1;
// music[3218] = 256'ha5d614e46ee267db10e32be25cd702d969db7cdde8e45ce675e971fb5303d3fa;
// music[3219] = 256'hcb02a10781002f067702d3fcd302600082ffb40486055f070b0e4b09d4fcb903;
// music[3220] = 256'hf7073b04130dcd0a72064711700a50fa4df956f24dea60f0a8f04bec6be8a1e8;
// music[3221] = 256'h02f5a5f9d7f4acf339f604ffe204a106aa09a50ad8075002f6faeff57ff9abff;
// music[3222] = 256'h17020dfd70f6abfff20399fdfa000e0179005008c30abd059306840d8f099203;
// music[3223] = 256'h36034401dd01ed053a122619a114f415ed10c40c0516e3176c14fb148c1ad721;
// music[3224] = 256'hc120bf1f5c2114204125182756256a30d1349b2fcc2be824a729ca2d272b4f33;
// music[3225] = 256'h5f33072e3732be371f42ce4c2a4c77471f4d8e4e3847b04b264d81461e47b147;
// music[3226] = 256'h3c47ef463847dd475a478844ae3ee241924b714e504a9944134143333023d421;
// music[3227] = 256'hbc266730c935cd2f5a2d022f342ffe2fbc325132202cab2ab22ebe2c1e24ce1c;
// music[3228] = 256'h511afb178916d9195316bc0bc8095507c8fe5efbe1fc4800c3fd4ffb29fda5f3;
// music[3229] = 256'h9fedf4ec36e47ce5dfe4e7dc1ae1dbe146dc9cd622cef0cd12d071d258d8e6d3;
// music[3230] = 256'h89cd60d033cff0c409c296cbf7cd7ecaf7caf5c8fdc737c785c806cb9dc23abf;
// music[3231] = 256'h9ac7c6c9c1c51cc1f2bd81bbfcbb58c358c3c1bc93cbeee221e2e5dcade0a7df;
// music[3232] = 256'h17de9adc7ddb41d6a7cfd1dbf3e2b1da42de89e429e302de13d81cdd3ce7f0e7;
// music[3233] = 256'h80e4bbe46ae421e4ddda5bca0dcd91d52ed404d2dfc859c459c6eec6a8cfb0d2;
// music[3234] = 256'h5bcd18cfafd1d1cf06d147d714da24db46d874d074d3f9d5fed26cd504d1e2cf;
// music[3235] = 256'h23dcc3e0cadbdbd685d2dcd3afdaaadba2dd87e2e6dc67db6bdf62dc33e115e9;
// music[3236] = 256'h62e227d300d20ddfc7dfd4df48e7cbe2b3e3aeef38efcae6b4e425e322dfbae1;
// music[3237] = 256'h5de1ebd425cd7fd6c3e2a6e3bfe5ceee2cf628f7d8ee59ece4ee0bed6bf0c6f0;
// music[3238] = 256'hcdef5ffc740b7b0fbe0ecf1201121811a712a90813082c110711e61212158e18;
// music[3239] = 256'hef1e8622a52953308636a4386a36fe3cf63f094005413f344f2ec331292d412e;
// music[3240] = 256'ha130b62fa034453546324337fa3ef23ba3386e3d1e39e939b841843de6416446;
// music[3241] = 256'h9540aa43ce411b3ca2429e4a9f4a1a4668434641ae4259453b45184669431f43;
// music[3242] = 256'h8f43543e973c93385f3a743fc935a334513a1d37883ee43e742e3f33073c462f;
// music[3243] = 256'hdf300d391f314c2ff92da02e0239e2367734ea3a90382131682d6430ab31872f;
// music[3244] = 256'h8830672b5e279927d221bb1e6b1872153f25bd29011e861a181ad21711156a13;
// music[3245] = 256'h33147613ce11fe09a104930a760302f4f1f59bfe57031d04d8fe52f8cbf1e7ef;
// music[3246] = 256'h9ef775f50de0c8d0e9ce60cf55d1d6cd20c71ec6c9c747c629bee9bf5bc9d8c8;
// music[3247] = 256'hf2cfb1d19cc46ec95dcb62c119c64fc7c3c28cc329c480c70ac23cbdd1c700c9;
// music[3248] = 256'h00c58ac66ac1d8bf93c2fec226c317bf0dbedabde0b95ebbdec070c796c7c3bf;
// music[3249] = 256'hddbe5ec187bf71be97c0cec3f1c3b1c3a9c521c597c5e5c93acf53d35cce21ca;
// music[3250] = 256'h42cf55ca31c3fec565cb1bd5b9d7b5d51ed1afc6a7cbbecd07cbffd358d515e4;
// music[3251] = 256'h28f67df0dbeea8e966e442e92fe6abede2f862f364ef58f361f7a4f405ee3eed;
// music[3252] = 256'hfaf15ff759f812f594efa8efe3f91a0172fe01f7dced63e5e4e5cbef25ed21e1;
// music[3253] = 256'h35e424e84ce25ae40ee2e5d235d7dbe755eb4af20cf866f703fb2df6aff751ff;
// music[3254] = 256'h13f8e4f6d1f8d5f322f07be90eea3fed9fede0f2e6f130f04df4eef722f9c3f8;
// music[3255] = 256'hd5ff2d046eff96fce7f959fcc8012a089813e31078035907441667189314a51b;
// music[3256] = 256'hac1f171d9320a0243126dc259329382e95258c26563549327b2b8130192c4d21;
// music[3257] = 256'h96272e3425330b31e13104369d48c552cf4db250be4f8848a74a0a4b574a1c4e;
// music[3258] = 256'h9c4aa048bc4c684c7e4b6e4a824846482b4c694e7c46f948fc4c1d463e4f7e4f;
// music[3259] = 256'hae3c5933f12cd92d1030c62ed02fb72abd2be7271d1e8e251f2941285d2c582a;
// music[3260] = 256'h62268a25dc291c2dd72bb025d51de71f691eb218ca1718132b16661c6d1a101c;
// music[3261] = 256'h9618740b880644089907b80a440c37072e075502fdf48eef50ef2aec73e7e0ec;
// music[3262] = 256'hf5f494ebace489e5fae4e6ec07e897db00e23ae361dd73dd0eda52d59bd179d6;
// music[3263] = 256'hfadb12d515d5e9d648d4a4d80ed37fca42ceb9cf94d0b3d052ce79d89de7eee9;
// music[3264] = 256'h6ce67de8f0ebc5eb5fe8e1e384e65fed69edadeaddeadfec76ec95e743e8b7ef;
// music[3265] = 256'h93efcded22f30df01eecd7f0f3e577d585d33ed40bd490d34fd828da55ce1ad0;
// music[3266] = 256'he1db3edbacd7f3cd99c2c3c799cfe9cceacd95d1a9d266da5ed985d182d8eed9;
// music[3267] = 256'h37cd99c74ece73d5b3d77dd8acd552d693d9f8d7d3d81bdbb4e07fe0f3d98ddc;
// music[3268] = 256'hefd709d354d948d598d028d8c7e034db31cf28cf91d3c8dc19e313df08e7dfed;
// music[3269] = 256'h36ecf0efede643dd21e153deb5df45dfdcd023d3abdb07d945e0a8eac5ee29f0;
// music[3270] = 256'h1af028f27def2ef1ec02910cdf02d1fea205e709d90c500b090a960b780312fd;
// music[3271] = 256'h66ff33078b0dbf07be0b5f177718ea1aa0184b185b1f571c721cb41db712c10d;
// music[3272] = 256'h54140e1ccb184a0fbf14551b1614c813ea1c8a1e141f2129412b4b243328a62b;
// music[3273] = 256'h7b2df23478322f2f133287368f3ba233902c0f2d38298d30a9385f336e2f5c2d;
// music[3274] = 256'ha131a33932377438813fee39a232942d802229290e362c2bcc277330192dc527;
// music[3275] = 256'h2b25152b1934cb31e62d352c4e2c51270f23c52998280227bd286b2654286b23;
// music[3276] = 256'hb226c42ce924ce295d280720c5239d1e861a821cb322fd2ec82f452a70273226;
// music[3277] = 256'h4820881cc620721dab196517ca123411390aa00419002e019c0739032203d402;
// music[3278] = 256'hb3fbd9fa9bfab2fc4ef4d8e1badae4d976da18d867d663d727d2b4d0d6d2fdcf;
// music[3279] = 256'ha6ce5fd21dd269c9c0c651cbbecb51cbf5d177d3accb3bce62cf92ca35cbd9c1;
// music[3280] = 256'h19bf98c4fac2e5c89fc99dc5a4c6c6c1f0bf80c2e4c6a5c523bf58c47fc5b4bb;
// music[3281] = 256'h09b948bebac129c042c1cbc103c357c8b3c56ac419ca14c8b5c3f3c740ccfdcc;
// music[3282] = 256'hb3cca4c8a1cb17d123d1d1d679d3b1d323e1d1de6dda0ada49d9d4dd76db30de;
// music[3283] = 256'h87e12ae71afabcfa53f52dfd3aff0701450365ff06fa31f860fbfdfe49ffaafc;
// music[3284] = 256'h3ffe6502fa06c50b76087b039801a4ffc3ff0d079e0cd7f80feab6f1d8ef8ef5;
// music[3285] = 256'h82f9d4eaabf4c8030dfce1f71af69df1f8f056f287ef96ddc5d7e6ecaff454f6;
// music[3286] = 256'h8f0055fc6cfe2d0948074405a602fb00470169fb64f8e7f855fc2cfddff712fb;
// music[3287] = 256'he7041007d2fdbbfcde082707befe68ffe9ff6302f508a50cf60ceb0c7509f109;
// music[3288] = 256'h800e3d0a13099a0dae11d519c11a59168e130417081fec1e23220b263823f323;
// music[3289] = 256'h54234f279a2be329432a322891299c2d64340042b344204056447f4b6c485c45;
// music[3290] = 256'hb94bb74a904aef4c124a674ece4ec84a6d4d0b4ff64bfa47bc4c054d1a452447;
// music[3291] = 256'h314d7049c23512282730fe3324312c32fe2ff829cb2895281a270e2c31286d20;
// music[3292] = 256'hf525d82610247625072807288e25f128762747261b26381bf11b261f321a8b1b;
// music[3293] = 256'h8115e60cff0ade064f07fa08b2003fff5406c601d2fc42f74bea66e998e991e3;
// music[3294] = 256'hcddf93dc2adea8df11df00dce0d7fcd7add340d41edb92d9a1d12ccd25d263d2;
// music[3295] = 256'hb9cad4c900cd83ce20ceaccfa9cb78c432c677c817ca5ec852c47ac27abe1fcc;
// music[3296] = 256'hd9e08ee107dee7dfa2de58d75cd71bdfd5e071e0cddc65d9c1d9c9d6c9d62fdb;
// music[3297] = 256'h09dd5cdb61dffde16ada33d81adb66e100e03bcc0ec5bdc6a5c38ec85dcceecb;
// music[3298] = 256'hcecbb1ca43caeacb30cc2bc6d5c6dbcbcfcc18cf44ce6fcedfcff2cfa0d3f7d6;
// music[3299] = 256'hc2d8e3d2cecee7d43dd65ed80bdb22d8bcd578d2f5d343dad9dedddeeddbf3db;
// music[3300] = 256'h0bd9d8d6e8d6a8d89ae037ddb4d6c3dbe2dc6bdd6bdd33dc4ede84da74d80ddb;
// music[3301] = 256'h24de05e546e662e43be542e787f068f4feea9de71fe994e4bce3dce523dda2d1;
// music[3302] = 256'hd9d679e0f3e167ebb4f0d8ee2400a80e1b0fd5130c10ee05cb065b0a9308160a;
// music[3303] = 256'h810a5d0033fdf601cb041a09a20aeb0a4908f209e4136e178b1f442573233e21;
// music[3304] = 256'hca0b7d04231a27218022b5260425d129b32f702df92a212cc52e76347237bc36;
// music[3305] = 256'ha238173ae23d0e42d83fc93a2b3c6a46cd457e44c24c4e444c3ea6460346f747;
// music[3306] = 256'ha14bc04501423941673f2242b54569459043484179453b46653bb63bc5404e40;
// music[3307] = 256'hb142413ed038603a3e3c873bef3bd04358452b43ec44413ec03d4d40c2361532;
// music[3308] = 256'h6033d134de372d390a3c8e3ddf39e538a8383334cc363936402f673bc0480846;
// music[3309] = 256'h78420e3e1a3c11396735d533f52ee130612b341f1421751fb61b6416450af509;
// music[3310] = 256'h490abb040b06bc066c02e101640145f207e0c9dafad8e0d558d538d7b3d58bd3;
// music[3311] = 256'hc0d5f7d412d16bcf57d0bacfcfcab7c804ccaaced4cb39cb39cb61c689c605c8;
// music[3312] = 256'h27c96bc73cc3abca7dcb39c90ecccac49ec479c3b8c27fcc95c235bceac51dc7;
// music[3313] = 256'h34c8d2c5a4c268c37ec0abc241c559c11ac0cfc40cc93cc612c254c264c34ec4;
// music[3314] = 256'hf9c6ddc594bf78c19fcc88cb5ec04bc22bc82dc69ac25cbfaac6abcd9fca7acc;
// music[3315] = 256'hf9cc10cc5fcaaac989dbe4e665e2c5e5e6e753e7b3e945ea3deccbead7e8f6eb;
// music[3316] = 256'h51ea83e98defacef32ee61f033ef7fed39ee86f3eef7c1f4c9f3d1ef8ae31ede;
// music[3317] = 256'h07dff9dc90dcfcdd66dceddad1dc03e441ebf1ed59f2fdf19bee63ea68e1cde6;
// music[3318] = 256'hbcebb9dd04d637da56e102e130e34cf409f947f88001c20035fb5cf979f4e5f1;
// music[3319] = 256'h80f6bef77cf2b9f028eed9ecb1f1a3f12cf02af57ff88df675f325f027f1c6f7;
// music[3320] = 256'h07fbb6fe2c034202b50177024806060e0113ea14b2161519ce16e8153f1c8a20;
// music[3321] = 256'he921b21ff1202229412b832ce6284923a92b582c962cd33fb94bc44d704d224c;
// music[3322] = 256'h3d4f844a254b1e53284c91483b4d9a50d3548553c1538551554b534d864ea54f;
// music[3323] = 256'h194ddb437b471e54a04f2f375029af286b245c26c82b3a3339352d2df2311d35;
// music[3324] = 256'h3e318532dc315432c12a4527672e5b2a252d4b33bd2e762d7731fa34142f312b;
// music[3325] = 256'hde2b6b2784292025aa1bc91a8818ce190616f40a290a1e0e651154120210630a;
// music[3326] = 256'hcf045108c207b501bd00c3f8daf2dff96cfc0ffac4f75ef165edc1eaabe551e9;
// music[3327] = 256'hf1eecbe884e603ea28e78ee4dcdc0ed8d6e188e2b7de23defed760dbe8de0fd9;
// music[3328] = 256'h74d573d79ce5f6edf1e635e70bedbfededed6feeb9e743e38ce63fe369e480eb;
// music[3329] = 256'hd5e687e16fe206e505e91aea3ae657e9f0ef4be9d7e9ceec27dc9bd514d75ed3;
// music[3330] = 256'h89d5b0d5dad710db54db04df73e154e1e9da1edadae1dbdd0bdb63dedcdcc0db;
// music[3331] = 256'h90dddfe168ddf2d2b6d280d23dd18fd6aed644d3b3d744d86fd1b6d0b4d195cf;
// music[3332] = 256'hc1cf18d244d5ded774daabd843d448d313d066d116d846d676d561ddece00cde;
// music[3333] = 256'h8fdf1ce03edb03dc36dd1cd9f9d776dd2ce4b4e296df57e168e645ed6eea2de5;
// music[3334] = 256'h5fe542e22be43ae95be01ad067ca65d06ddeddf26dfddbfea104480a240b9f06;
// music[3335] = 256'h29078e0bed041a0218067005fe056f04b901f702ca028f06020b5105ad025e08;
// music[3336] = 256'h260dd011240da00150fe38fd48fd2403c209120ba20c2112480f4e0d0d11b413;
// music[3337] = 256'h101970157818f323d21df61bf1209d22ce29212a21276229172d8e2d4f2d9430;
// music[3338] = 256'hd42b2d27d82ed533072f0a2cc730e5309b2ff62e672e3235c9347a35163a0f31;
// music[3339] = 256'hfd2d0c2f4d2e0934a9335131af334534fc31ba30f8312b31002d522bfa349835;
// music[3340] = 256'he229c32eb62fc825c728662edc2a3126442a942cc42e4932052a142bdb2b382b;
// music[3341] = 256'hfc3e2e43143de940c23b05372d320c2fa4334132fa2d222baf22881b261f711e;
// music[3342] = 256'h99167016431447110c10820c0410c112cc0cecfcc1ea28e71ce9f8e65ae120dc;
// music[3343] = 256'h1dde5fe111e20cdf55d9c7d54ad5c5d641d754d791d285cda7d2c9d285cb2dc9;
// music[3344] = 256'hf8cc06d437d2eacac9cb7cd04acfdac605c69fcadfc739c91fcb69c825cafcc8;
// music[3345] = 256'ha0c9a7c985c04ac399c734c1fec433c586bec3c178c33ac6c5cb43c771c396c4;
// music[3346] = 256'he8c134c33cc87cc758c958caf2c48cc707ca7ec51ec544c762c9b1c6a6c6e9cc;
// music[3347] = 256'hfaca33cc49cf41cd33d2f0cf09d44feff9fb02f7ebf78cfa79f83ef712ffeb01;
// music[3348] = 256'h62fbdcfce7fce9fb100206fea2faeb004700960000ff20faf7ff8d0065fff704;
// music[3349] = 256'hfafb77ed4be7bce737edcef0f2f5f7f2ece5c8e65aede2eaf8ec2df425f456f6;
// music[3350] = 256'h5f007204fd03c6fd7cf461f690fa83f536e536de4eec81ef66f09afe15045a05;
// music[3351] = 256'hee088809440948086e04570115067b0586fd09f855f646fd67ffe0fb59fc8afc;
// music[3352] = 256'he60103048503df09700d7e0d970c33101015a016e617ce15bc16a1154212e812;
// music[3353] = 256'hc20dd40dc413111a881e351d9620a920fb2054220f209828f924b62a1f45bb41;
// music[3354] = 256'hc33ce54434446744e44125497d4e1144d6459d4aa8467a458a4569448d458b49;
// music[3355] = 256'hfe496f49704c7f4c6f47e246224a343bf6284e2cee2d7a2c73349e324e2d5130;
// music[3356] = 256'h0e2d832dc936e43374314f355430b22f0332cb2d232e4f2ee02a8a2ab22c5d30;
// music[3357] = 256'he8316331e3318c2da1265822332094247523b21a281f2023db1d6a1a5b12020f;
// music[3358] = 256'h8c102d0913046203bfff06fd20fea6fbb7f277f191f6c4f373eed2edeae94fe2;
// music[3359] = 256'hede2cfe419de68db60dfa7ddb2d4b5ce65cfd2cf6dcfead061d184ce9dcae9c9;
// music[3360] = 256'h25ca6dca36ccdbc8c1c82ad76ee019df03e151df17d9a3d712dd1fe1bbdb52db;
// music[3361] = 256'h0fda49cf57d3f2dba1da67dcdfdabad8c9da32da4fdb90dafad9b3dcbed0f9c0;
// music[3362] = 256'h41c29cc3d9c30dca29c65cc32bca80c927c735c88ec85acd12d07ccabdc9ead2;
// music[3363] = 256'hb6d300ce8bd2d8d297cda7d08ecf16d08bd82ad773d523d7efd0a0d087d492d3;
// music[3364] = 256'h1bd540d847dce4dc22d7f8d294d329d521d171d183d8aed7e9d6fbd82edbabe0;
// music[3365] = 256'h60e1eee052e31fe5c4e2f1dcc3de73de68d94be0eee8fae4b6dfbae293e27fe1;
// music[3366] = 256'hf5e5e3e3cde60af0caf141f293ee7eeb82eb8de43cdeaddb57e243f1ebf6b8fa;
// music[3367] = 256'h3607f50e090e330e3c0fb911ca14d90d9d07b90a0f0aff08460a990587046c0b;
// music[3368] = 256'hdd0dfe0b520922093c0a15ff47f603fae5faa3fed9023c058505f8008709390e;
// music[3369] = 256'hbf0b921a072255201f259f2a5731753390339b33d9322035ef35e839493bf738;
// music[3370] = 256'hfb3b393d3d3d443c193d2f42e63e8c3cfb44d5477e4399450b45d7408e478446;
// music[3371] = 256'h273fdd447d4550420247f348bc456942f2439644fa40ff3fb140e63f163eda3f;
// music[3372] = 256'h5443493f81377a3470398f3fba3c033b583f4f393c32d7342837da3c393ead3c;
// music[3373] = 256'h1f3ff8372a4207568a535556a955544ecf539952ec50124de644df44da3daf3b;
// music[3374] = 256'h873f1437a934003a4238d032af2dde2347172f121814d912540146eee2ef80f3;
// music[3375] = 256'h0aec93e417e343e394dda9d9eada51db1dddcede0bdde5dd9edff6da4adaacdd;
// music[3376] = 256'hd6da05da2dd7add20cd4d4d00bcfa8d095cddfcdb5cf18d0b1ceacca76cb6acc;
// music[3377] = 256'hc0c88fc4a8c03ac26ec757ca75ca73c50ec2c6c078bbb7bdd0c578c7fbc311c0;
// music[3378] = 256'h03c126c056bbeebd8fc467c4a3c0cdc614c9e3bfcdc147c467c377c690c5c3c9;
// music[3379] = 256'h6cc758c260c900c9aac987cab6c5c2c7f4c800d670e98fe9ede567e5cde2f5e1;
// music[3380] = 256'ha1e4a6e746e8c2e8f7e66fe498e2ede242e915eef2edd4e9f1e97eece8e901ef;
// music[3381] = 256'h91f1e3ee57ed9cdd35d6bddbabd915db04dbaed8e5daf5de77e3f2df32dddadc;
// music[3382] = 256'h83d82ddc67e059dfeae3b2ed2ff47df646f4e5e917e6f2e6bce1c7e5b6e13dd2;
// music[3383] = 256'h31d609dd03dd6ae4a8ec7ff313f878f7b5f6dcf512f338f3f8f6a1f638f44ff1;
// music[3384] = 256'h47eba5eadceb9fe93cee47f299ee34f155f9e8fafcf9a7fcbc005e05d4042e03;
// music[3385] = 256'h2d0b120d310c44156c10220b2b17361b971a121b3e1d9922071fac239c2ad224;
// music[3386] = 256'h6d30b043d3461c44c3400740294289455f48c045b9410f45384e324f7a4de650;
// music[3387] = 256'h0c4d5346d344e447e74ed250f54d904c3b4d0d4cf540fe34dc36ea374331f035;
// music[3388] = 256'h8b3877300c313a33b435da34ac2c7835323f57386933c635233a9e34c42dd031;
// music[3389] = 256'ha631672d5e2eba31bd2d2c28c12a172ef231ca30c32a2128ab225e2064208121;
// music[3390] = 256'hf922911b8919a5199a159516f312350e150cee0662026105620e9e095b026e07;
// music[3391] = 256'h21073304890576024af9edf392f502f593f41bf213ef92f07bf03bed72e765ea;
// music[3392] = 256'hdbec5ae198de05e1d1e077df8ee061f15bf7eef153f582f407f695f4ddee86f0;
// music[3393] = 256'h83ee7bee6fefe9ecd2ecc2eac9e8d9e989ed42eb70e546ea9bece4e700e463e4;
// music[3394] = 256'h32e5ffd7a7cc4bd155d586d495d21bd3bfd70edbb5d7e8d31dd8c5da13d74cd5;
// music[3395] = 256'h30d59ad33ad5cbdc9cdfd7dc06ddedddf1dd8adb61daa7de06dd44da82dfcadd;
// music[3396] = 256'h29dadadbc5d3a1cf50d4d7d2f2d349d37ecff9d0e1d34ad95fd595cd95d054d1;
// music[3397] = 256'hc3d0c4d31ad735d6b5d4abdaabdab4d96bdcadd8ffda45dc69d86bdcf9e0c7e1;
// music[3398] = 256'hd2e093dce4d6e7d839de16dd58e34ee8c7e4cee752ea3eee6eef62e958f328ff;
// music[3399] = 256'h9cff78fe44eed7e18aee6bf840f91c00c50adb0d70089608e10ac309db0ade08;
// music[3400] = 256'h9706fa04cc03dc04a101b402c304a0fb7df1a4ecc5edb3eeebeeaff494f969fb;
// music[3401] = 256'hc6fcee011c056103fe089e0d27100912a90df9115615d613621b451eea1db922;
// music[3402] = 256'hec258d25db22e421542296262b28832145229c27d22cc334eb31cd2c06312534;
// music[3403] = 256'hc633e433f436a7363d322c33973238318e32472e062d113041327e36a833e32e;
// music[3404] = 256'h1730c72de82ba52f1433ac33fc30ee2eca2f222c4928b6309736662e452b0032;
// music[3405] = 256'h5730cd29542c772a3629ce3af84547455a48bd47c747a048ce435c41fe43dc43;
// music[3406] = 256'h1d3dd23b523c84357e339c32472c3c2a282b11272224ab22aa1ac31a29179d00;
// music[3407] = 256'h11fa0afde4f427f3fff2e8ee13f09cf2f7eb89e4e5e67be448e2f1e4a6e3f7e2;
// music[3408] = 256'h6ededaddf2df1eda5eda49d702d260d542d6e0d7f1d382cde1ce7ccafac629cc;
// music[3409] = 256'h91d06cce33cb4fcee4cddccb6eca2dc81acd38cb73c74dcc14c721c357c75bc3;
// music[3410] = 256'h5bbff9c21cc62ec415c39ac691c742c67dc680c7aec9ecc807c4e4c17ec459c8;
// music[3411] = 256'h7cc842c50fc334c222c420c705c964cbbbcb26c9e8c3bccaf1e044eafde828e7;
// music[3412] = 256'ha4e171e5cee829e6a8e772e954f0e6f71bf9b2f7aef53efa1afe14f919f8b4fd;
// music[3413] = 256'hfafb55f831fee6fe64fbebf646e835e137e6cdeaf9ebeeea89eee0ee5aefbaf1;
// music[3414] = 256'h8fedcdf203f7ebf195f33ded11e83bf3f4f755f7f9fb87fdf0fe74079e0d5a07;
// music[3415] = 256'h0301e2fe1ef6d6f5a5fa34e92adc4de664eecef558ff3d032c068c077008fd08;
// music[3416] = 256'h850728070904d4feefff3d02dafc9ef742f8a9f8d3f92bff5602d8fe49ffe105;
// music[3417] = 256'had067106a70a350ef50e650f7f13c51429140318261bf61c8f195e15e1167a16;
// music[3418] = 256'h09175c17c21a362aa23595378138ef3a603e7d3e2f3f1d3f873e4e445745a841;
// music[3419] = 256'h2b42b6420247064bbe463f45af487f4a134c664b744ced4ff5451a367436dc3c;
// music[3420] = 256'h013ad035d93612363a327b34463a0d3a3f36e8330a34aa33452f832c1b315138;
// music[3421] = 256'h1d382132c7313b31432c2a2b052ac128682710247c276f294b27042a232a9f2a;
// music[3422] = 256'h9b2b75262b24c225ad269323671f751f5d1bcd169516b91370129610590a3d06;
// music[3423] = 256'h0d0471ff4bfa6bfa01fa04f40ef34cf4c8eddee7afe5f3e3f6e686e56bdd18dd;
// music[3424] = 256'hecdc70d95ed94fd8efd892d67bd2c0d359cfd0d130e142e5d8e077e0b2e2b3e3;
// music[3425] = 256'h5ee0f5de79df07dd37db0fdb0fdd3ddfbedd7ddd84dddbdaf1d8b4d7e2d922db;
// music[3426] = 256'hd0d728da53da12d075c674c268c3cec424c5bfc7c4c7dec485c609caf1c612c6;
// music[3427] = 256'h4dcba2c8d1c4afc896cb82ccf1cb30ca2fcbf6cd6ace30ceb3d0a5cfb9cb12cb;
// music[3428] = 256'hddc970cbaad095cf25cc57cc9acdc5d094cf72cd33d4e8d424d35fd79dd33bd4;
// music[3429] = 256'ha7d896d2a8d20ed7c7d6f7d53fd39fd211d3f5d386d8ced88dd696d877d856d6;
// music[3430] = 256'hb4d8badac4da37dc2ade16e03ce153e083db57d83edd6de0eee0d7e51ae67be3;
// music[3431] = 256'hf4f2b70af90d2c079f04030091ffbe00d1f854ee2aede3f435fe44066909dc0a;
// music[3432] = 256'h6a0e97101d12c710dd0f370fa50c9a0ce00af60a22059bf6a3f232f0ceee62f3;
// music[3433] = 256'h1ef357f56ff6f8f6fcfcc4ff3b00200136061308b404710a490dca0cf611d914;
// music[3434] = 256'ha61c56270b2a8d2ad82b8e2c052e8d30be306b32d6371f39b03a013fe83d0e3d;
// music[3435] = 256'h9f3fc33f1641ac44d043d33f7e3f94418342db441a4635445d447a45a5441c43;
// music[3436] = 256'ha244b0483f475f44364543458f432d405c3eb9403446d1485244ad43bb43983c;
// music[3437] = 256'h0739d93e8349ff48ed415742cb3ddd42ba53fa54a6554a57aa52a1568c566052;
// music[3438] = 256'h20542953eb51f04ea64d6750d64bf548c249b445c8426b3eb939923a643aff39;
// music[3439] = 256'h5e375e284a1ac917af127a103912380593f934f9cff371ee9deb12e920ea27e8;
// music[3440] = 256'h2de5b6e5aae354e072e13be39be1c6df10dcc9d625d59cd3acd248d327d137d0;
// music[3441] = 256'h72d0becfbfcd59c866c754c97ac6fcc5b3c63dc517c774c9a4c64ac49cc5ddc1;
// music[3442] = 256'hc4bfbcc480c3d8c108c3f3c19cc249be18bb3fbf91bf4cbf20c005bf74be82be;
// music[3443] = 256'h27c13cc304c29ec179c20bc2efc130c2eac291c636c778c605c699c365d289e5;
// music[3444] = 256'h81e542e64be75de3b9e3b3e0c7e1ebe734e782e75ee995e88be9fee727e4a7e5;
// music[3445] = 256'h7be81fe985e8f3e6aeea16ef5bf020ef1ce1a2d552d81dd740d5acd7c7d795d9;
// music[3446] = 256'h82dc26db3fd722d95cdb21d8ecdb92e03cdd84dff5e5d8e3eadcd8db62de35e0;
// music[3447] = 256'hc6e379e4bbe298e64deeeaef49e9e9e47ee1a9df3ae5d7ddeecdbbd013db57e0;
// music[3448] = 256'ha8e6a9eefbf319f55ff501f60efafffaf5f3bff2d1f2cbef77f175f07cef9ef0;
// music[3449] = 256'h0fef1af1a3f2adf1c2f3f8f7fefac9f87ff9dcff070048ff27038f037204150a;
// music[3450] = 256'h8c0b450c6d126112d81262226e2f3833c037043786343b37b639133c7d3c3e3b;
// music[3451] = 256'h063e44412e429a42a5443a48694739443646a14aa14cdc4b2d497b4a9a4b4740;
// music[3452] = 256'h6f37d73a5239f737663ce23bfd3bc13d043b9137ee356c34633160330e3b953a;
// music[3453] = 256'h2e352e373038ea31a42f85350d3a6d37673349317b2d712c5c2ed62d042fc52e;
// music[3454] = 256'h7f2cdc2f8831e62de92ccd2da32dfe2b9e271525f826f225df21be1f8d1e171e;
// music[3455] = 256'hee1b671584101910720db707c80223fee0fc0afdc1fe16059605a6030a0453fe;
// music[3456] = 256'he1fbbbfe1ffc38f74ef7acf6b6f028ede1ea25ec99edfde901f679010dfd24ff;
// music[3457] = 256'h09fef8fa70fd7bf9fbf62cf524f213f305f3e2f27ef159efc5f169f432efbeec;
// music[3458] = 256'h7bf284f113ee1aee6bef71ee88dfa9d573d9bcd9f8d796d5f7d5c7d809d9f5d7;
// music[3459] = 256'h46d3e0d367d6fad496d83fda40d840da14dde1da23d85bdaa4d8ebd620d8c3d5;
// music[3460] = 256'hadd6d2d7e3d9a9dd9cda5bdaefdc7cdc80ddd5de6ce3c0e5c9e25ae3a8e1eddf;
// music[3461] = 256'h21e1cad87fd098cfbccf13d3c8d0ffcc0dd187cf75ce6ed441d675d272ceb7d1;
// music[3462] = 256'h06d6b8d40dd406d4ead67ad955d860d913db19db36da96d9d2d99add73df51d6;
// music[3463] = 256'h19d59ddae9db0aedfafa9cf76efe1f07190541013ffed3fb8ef8c3f915fa75ee;
// music[3464] = 256'h2be7d6ec07f3a2face004302f3089b0c9a0a420d350c3f09a9033cf49eec30ee;
// music[3465] = 256'h94ece1ecefed7dec02ec03ef91f3dcf335f3c7f503f8c2fb0efef8fe8f057006;
// music[3466] = 256'hf6032009f807bc07ae0fb7118312b7146e17a9199b17741afb1e162141235822;
// music[3467] = 256'h9c24a126f8243326b22724280c2720284d2b8c294e288529a42db331ad2d922b;
// music[3468] = 256'h482fab317c315c2fd730c831b82ef12ef1310f35d3349d3187304d2f5d2ef72f;
// music[3469] = 256'hb532b232e12df62d2832b22c2e25bd27642ca234dc432e4a59484f4735436a41;
// music[3470] = 256'hb042e34315460946a745d744db449f47b5457e41e440d6434547f6441c3f173c;
// music[3471] = 256'h0d3bc13908394032de2109164d149713cc0f120d900ada035fffb2fdcdfd3bfe;
// music[3472] = 256'ha4f92ff9f6f706f2b9f084ec1bea60ea31e699e3a2e16ee0fddd03dc74db82d5;
// music[3473] = 256'ha2d565d8f5d58ed4cfd018cfc0cfbdcd5dcde4cde9cd51cd46cda9cbefca93cc;
// music[3474] = 256'h96cb51cc66cc0cca7fc89dc5d4c6a6c7f9c53ec81bca02c9d4c6c4c5e7c2dac1;
// music[3475] = 256'h08c681c56dc4d5c6abc898ca39cbd5c92ac774c8f4c72dc679c841c50ec73fcb;
// music[3476] = 256'h9acd17de50e52ce193e4c7e40be384e464e680e536e658ead4e7c5e71de8cbe3;
// music[3477] = 256'hcee572e80bea7ae953e986f6ab0088fbd5f9880198fd73eb3ae3f3e51ae8a8eb;
// music[3478] = 256'h31eed8ed1dee31eef1eee9f01bf275f4c1f24cef32f220f1a9ee45f0f5ef5af1;
// music[3479] = 256'hd4f242f47af193ec4df239f4d7f381f97ef8aaf82cffc304ae022bfbbdf91df6;
// music[3480] = 256'h99f3cef5acead5dd26e496ed27ee5cf65e0076ff5002c60478033705ed030a02;
// music[3481] = 256'h8502b503fdfe23f90afdf4fcb4fae1fb38fb67fdcdfe1b029404f603c007100a;
// music[3482] = 256'ha90d2a0f6c0f2214de128a16e9197c1cd42ee1386d38b837d32fe52cb02f3334;
// music[3483] = 256'hd034d432433a303cd0374e3cf83e393e2b4291441a442445e245bd485949d847;
// music[3484] = 256'h454ce5440d34d72f5f307630d7309e33bb375f331e321d378c38b139913a753a;
// music[3485] = 256'h5439fa34ad2f2c3216396036183477332c2ed92dff2c0c30ee37f534ca315d32;
// music[3486] = 256'h2e31f62e6d284c27022b132964265025c7241e28bc2c1d2cba295d283f27cf29;
// music[3487] = 256'hd027cd23a925e421111eba1e111aa4144e104a104710b6071d06590792006700;
// music[3488] = 256'hb3ffbbf970fa83f843f334f1bfeddaeb4ce9b2e636e5e2df7edfdfde71de4eeb;
// music[3489] = 256'hacf0bbeb49ec3cea8de7c5e7cae790e79ce5cbe5e0e682e6f9e584e494e587e5;
// music[3490] = 256'h2ae09ddcc3dbc5dbf3dfdbe01fe0a7e375d9fec77cc414c57ac602c774c4adc7;
// music[3491] = 256'h9bcbb0ccf8cc50cb34c977c6a2c714cacbc638c4aec750ca1ac948ca5dcb42c9;
// music[3492] = 256'h31c976cacdcb74cb54cafaccffcea2cfedd134cfb9c742c613ca26caf8c7b4c9;
// music[3493] = 256'hdacd42d074d1c7cfc7cebdd203d1d6cd67d234d331d133d32ad66ed6fad288d3;
// music[3494] = 256'hb1d6e6d303d2c2d528d5d4d200d89bd91dd705d96bd9a0d9c9d8c3d8eddc47dc;
// music[3495] = 256'h81dd80e10fe07ae090df12e281f19afb56faf5fa50fede00b9016c06970f0d0e;
// music[3496] = 256'hb70501046d001affa90545ffbeed56ec35f923013d046a09310dab0fbd13bd0b;
// music[3497] = 256'hcdf9b4f6f1f787f3c1f443f2c1f0cdf48af437f7d0f6d2f34af648f5f2f5b5f7;
// music[3498] = 256'h70f765fcb9fd43fc27018b045803d0053f083b08fb0f5d14e1118b17e119d81b;
// music[3499] = 256'hd627d92b192acd2c1830af3298331136b837b438bf3c9f3b463ad63d7c3e6d3e;
// music[3500] = 256'h3e3f2c4092406a407c4330460d466e444f42b3437546fc460b47b34769479d47;
// music[3501] = 256'h18463b429c4398449943a7458c45e948dd488b419b405740bc457c503656cd5f;
// music[3502] = 256'h5c621b5d805b5c568255895620539c546c54c153ff571c59c359d257ed52ef54;
// music[3503] = 256'h4f53894e5f52864fc34bb54f9942812f072c1c28fb236826c9234c1f0b1e901b;
// music[3504] = 256'h001b5918b311b30cab09f10988010ef30ff09bebf5e891ecc5e7dbe689e5b7dd;
// music[3505] = 256'hd9de7fdecbd911daf3daf8d8ded406d28bcfa9ce4acc03c71cc9c4ca11c831c7;
// music[3506] = 256'ha0c4ecc59fc580c172c3b3c319c3a7c4f1c19ac07cc302c4c5c09fc1bbc272bd;
// music[3507] = 256'h09bcf1bcc0bc40c009c1cfbe14bf68c073c0c7c185c6e8c8f3c76cc6d5c4edc2;
// music[3508] = 256'h95c20ac393c065c9d7db62e10ee2d4e164dd2fdf0be4c4e527e596e551e428e2;
// music[3509] = 256'hade722e99fe635e8d9e637e852eaade9f6e9e7e6cfe637eb57e907dc15cfe0cf;
// music[3510] = 256'h77d30cd54fd7aad624d6cad610d881d8d2d8d2d9f5d771d9a9dc9bdafed697d6;
// music[3511] = 256'h6bd8c4d7ded950dc1fd824da08e17be2c2dfd4dad2da11e0b6e089df29e36ce3;
// music[3512] = 256'hcde4a7edb2ea69e30be69ee4b6e240e48cdf5dd37bcd90d6f2dd25e355ec41f2;
// music[3513] = 256'hcbf755f6c6f0f8f0cdf032f18eef96ebb6eb1fee2af2c6f188ef0df373f4a2f1;
// music[3514] = 256'hb9f08ef449f978f845f9f1fc78fbe4fd33039202f80cfd1e1f24f0239f23cb23;
// music[3515] = 256'he327d529812c0d31dd2ff12d9333963a253c143c2b3ce43b413dca40fb43ec46;
// music[3516] = 256'h3e4a3a484a487e48323aa232c237a1375537ce37233b773ca236653ac83d9c3a;
// music[3517] = 256'ha63db03d303da33f683c183be73bbf390037a9337936663b74365d332c34942e;
// music[3518] = 256'hc72a292ce430ae35f733d2315630152d912ace29322b1828e725bb2a502be228;
// music[3519] = 256'h5227a7269628a6284329242971252b244c234d21f4204e20941c681598108d10;
// music[3520] = 256'haf0f1d0db70adc06dc05060764028dfef7fc65f9b7fd90040504e9011cff92fb;
// music[3521] = 256'h2bfc5f04ba0d0f0e160b750900075a071006050099ff5c011bfec9fd3dfd7cf9;
// music[3522] = 256'h0cfaaefc88fd83fa3cf8d9f874f556f32df41df86cf6d5e234d80bdc09d93fd6;
// music[3523] = 256'h43d5c2d6efd851d753d9acd71ed4bed550d6ead80fd988d5e4d4add347d4f5d6;
// music[3524] = 256'h89d618d5d3d3eed5b0db43da35d489d309d51fd885d722d471d89eda18dabadb;
// music[3525] = 256'he5da65dcacd9a8d41cd82ddb61da36d880d7b2d8dbd892d9d8daf3dc3cdeb2de;
// music[3526] = 256'hfbdab9cf53cbd8cc0fcccbcd39cebacde6d1d7d32ecf8cd0cad63ad475d41ad6;
// music[3527] = 256'ha1d3e4d767d971d75ed9e7daa7d904d92ee6a7f335f53bf76cf26aec26f1c3f5;
// music[3528] = 256'h0ef87af930f8d2fa29064d0a0b027d016903edfdb5fc26fdc9f345eb55eeedf3;
// music[3529] = 256'ha9fdc602d4f682f343f8d8f6d0f900fbbaf815f990f825f707f43cf1b2eeb2ec;
// music[3530] = 256'hb8ed5ff2d6f507f211f27af7cdf838fa90fa4afc6f01e101b9ff51017606a209;
// music[3531] = 256'h540a700bb70dfe112e144215b9144412b917051d291b411d531f071c3b1c451f;
// music[3532] = 256'h33217724e025bb241e243a25b0287f29462b3b2c3127882a87303e2dbd2ce22f;
// music[3533] = 256'h0c31c630a03060308d319335d6357f34fa35db356c31352c0030df327432ef40;
// music[3534] = 256'hf94cbb482e474747e6442e4c69522e4b46496b4b3146b7474b4bc546c143f745;
// music[3535] = 256'h5d471b44b642e8439744a6451545d247de449734162a1a28602483216620311e;
// music[3536] = 256'h3b1c241b6d174e146910ca094b0aa30b10073c07fb05fffdc9faf4f8b9f421f5;
// music[3537] = 256'h33f3f9ed71ec03eb26e948e628e4cae29fddbbdcb7dcc5d7e2d6e5d733d71cd4;
// music[3538] = 256'he3cec6cd51ce4acbb1c7bac8b0cad9ca1fcd3ecc64c9aacad1c848c61bca01ca;
// music[3539] = 256'h8ec39bc21bc7c2c910c7dfc326c618c69fc58bc7c8c5a0c678c6e1c453c74ec5;
// music[3540] = 256'h5ac479c370c146c656c555c68ad5a3de7eddebdc2dddbbded5e1b2e01adeadde;
// music[3541] = 256'hbadee5e180e46be375e6b9e764e927eebeed64ecc6eb4aed80ee1eee0ef5e8ef;
// music[3542] = 256'h30dc22da84dd6dd7efdd02eb1beda2ed74eee8ec43ef71f00cee5def34f04eed;
// music[3543] = 256'h3deea4f0d6efcaf24cf42ff043ef7eedb0ec20f0eceee8edf1ef6df45af8edf0;
// music[3544] = 256'hf8eb12f23ef4d9f22df3b2f4bcf56af8020058ff24f77df689f4b8f152f7a6ef;
// music[3545] = 256'hdedd8ee29cedbded79f53dfe4600bb028f03a306c607e903a60333033c0013fd;
// music[3546] = 256'h5ffce8fe48fe88fdf2fed8fdc3fd6c000700ab02280b94088c07381962249326;
// music[3547] = 256'h172dba300432c73204330d359c38c73da741ee432844a63ffb396f3ae03afa37;
// music[3548] = 256'hb73bc43fa442d4465f448046424565355f2e7f32353365318b327934fb33ae33;
// music[3549] = 256'h0434ee36fc33492e2c330d32842d313157322d337533f3332e351230be2cbd2c;
// music[3550] = 256'h362e37327f32a131dd327c313b2d06296f2ad3319531412ced2c3a2996281b2c;
// music[3551] = 256'h0126a4259929fc28252a35298e2a902cad2cad2c0a2a5c2941261524c825a122;
// music[3552] = 256'hc820731e3e1a26166a0fbb0ee20e020ae009a60a7006290566036ffcabfc62fb;
// music[3553] = 256'hd0f3d1f2f1edc8f07b01f905010275fd0cfa62fa1df8b6f6e0f2d6ee2df1e5f1;
// music[3554] = 256'hebf142f023eb54eb2deba6e50ee609e931e694e8f0eb69e9e4e764db23ca95c8;
// music[3555] = 256'hbcca24c9b3c7f9c598c8a0ca08c708c8e4ca0ec6bbc3e8c447c240c32fc6fac5;
// music[3556] = 256'h04c530c45bc659c62ec21cc2cdc3a6c344c4b2c475c5d3c60cc6a0c5fbc5dfc3;
// music[3557] = 256'hfac25ac3f9c3cbc5cac4ccc2acc228c4fdc5e7c468c5b0c599c27dc31bc6b4c6;
// music[3558] = 256'hf9c8b4cae1c783c682c958c93ecb4acf22cd7ccd24d03dd160d308d305d40ad6;
// music[3559] = 256'h2dd62cd757d708d813d94fda58da32d952dbe7da53df3ceee5f3a4f2c6f4f3f4;
// music[3560] = 256'hf8f67dfbc9f80ef1eaf160f832faa9fd3100f4fd9e023909f5064203e3018800;
// music[3561] = 256'h9501e601b1fb89ef7be465e2b5e60aec4af13df59ef806fb23fdb1fd0cfc74fb;
// music[3562] = 256'hfaf762f49ff4faf229f2b1f1d1f0a4f092ed04eeecf0d5f02ef4b5f98efd4a00;
// music[3563] = 256'h5e0168027504810563072b0bab0ca80dd00f3512c3138f12df14b116bc192528;
// music[3564] = 256'h9930ca2f2e3190320635ef347d36103ac5361637053bc53b643d5b3f9b418a43;
// music[3565] = 256'h9b43fe425844b3468746b8460546e64476463c473347a4470f48e34713488a46;
// music[3566] = 256'hb242e6496c56035a935ba55ac758d659f156ee53ee51db51e7585b5ba5571a58;
// music[3567] = 256'h4057b2544954d2521954d656d457ec591a59f659395ca650134250406d405f3e;
// music[3568] = 256'h9d3e4f3c98370934d430ce2d362b6529e5251122b01fe91ae918c716ae0f310d;
// music[3569] = 256'he50ae907040808054303a3fb37ec35e654e587e25ae03fddbfdb11db60d80cd5;
// music[3570] = 256'h63d24dd17dd0e6cd1dcc1ccc3fcb6bcb32cb64c83cc867c8c8c515c4ddc2cec1;
// music[3571] = 256'h29c027be7fbf14c084be55c0bac1bfc0bec1e4c167c17bc224c20bc23bc2fbc1;
// music[3572] = 256'hcbc370c320c3b4c4e9c093c008c30ebf90c6ead490d731d9bbda67da56dc02db;
// music[3573] = 256'h1bdafcdad0db0ade28deacdecde1b7e4c8e5c8e3a0e348e758e80ee853eaece7;
// music[3574] = 256'h65e6a2e93bdf5dd191d234d4c3d13ed238d47dd4b0d262d321d548d55dd410d2;
// music[3575] = 256'h38d26ed30bd3f0d26cd0bccd4dcf88d0c4d03ed291d483d75cd7fcd5d1d6cbd7;
// music[3576] = 256'hdfd9ecd956d85fdafdddb1dd38d64ad4c2da0cdc8bdf93e4b3e23be5d1eb6eec;
// music[3577] = 256'hd1e73de46ae2f3df67e032dd66d001cc68d58fdad2ddfae62decf8ef2bf387f1;
// music[3578] = 256'hbef268f362f1e1f096efc4ef06ef40ec8ceb9fedf7ef6dee15efc6f02ef05ffb;
// music[3579] = 256'h8e0a980e2f1021132c15ae16c818141dfc1ef01ff4226023e625672be52b002c;
// music[3580] = 256'hbe2f1c359e398639c03ac83d7e3d7c40b241be37d62ed52e01307a30e331a331;
// music[3581] = 256'h2c310d320f3228330336a536603439332a34f433bf34da3530342a343f349635;
// music[3582] = 256'he339d13742360a3951352a32f233a93575369d331a31a930bb2e3b2c3a2bfa30;
// music[3583] = 256'h9a375035a531e02f9a2c182b2e297526b227bd2734262828ab2732253a264c28;
// music[3584] = 256'h03286125ea2541270e25f4247225cf236c21dd1f3a1f601baa18ac172415da12;
// music[3585] = 256'h870f2f0d1109010641059fff2d07e9127f0db0103c1af5167d140f15b1122f0f;
// music[3586] = 256'hcc0b410995078c066c05d0048005fd04ea01af00ceffbdfd8cfe50fbc7f9c5fa;
// music[3587] = 256'h5cec6ce0d8e10ae0c4defadf65e08cdf7fdd16ddf4da22dbbedcd9d9d0d799d6;
// music[3588] = 256'h4fd5e7d4b4d3dad2d7d349d65ad522d49ed4d3d2bbd443d775d501d673d63dd5;
// music[3589] = 256'hc6d591d578d447d555d619d649d6d3d64ad757d6d3d33fd35ed38ad333d58cd4;
// music[3590] = 256'h84d2c1d43ed72cd6f0d6b2d747d895da97d885d95ade1fde86debcde9cdfcae0;
// music[3591] = 256'h08d89ecf68d13fd317d2e7d375d5b2d3f6d3c0d301d4fcd3d5d3c5e01ceecfed;
// music[3592] = 256'h83ec4eed36eff4efa5ef71f28ef369f451f56cef73ebf5f183f788f9abfd7afd;
// music[3593] = 256'hbeff2307b208d4053401e801c6fedeef62e84fde92d3dadb8fe2cae6baefd4f2;
// music[3594] = 256'h66f76cfa71f82dfaa5fa39f7b2f1f5ed98ef67ede5e9b1ecd4ecc6eb40edc5eb;
// music[3595] = 256'he4eb4eef52f1fff2e0f5bbf8fcfa7cfdcdfd96fee4022a049203c005ef07cb0a;
// music[3596] = 256'h0d0fd1101a1181145b161215d116171afd1cc11e071f6220ad20af2187241725;
// music[3597] = 256'hff25dc288c2b572d462dc72cf92dae2fdb2f2e3117345034ee34b6364b366036;
// music[3598] = 256'hfb356e368e371a38a742014d194a244996496146d448174db54c864a4e48dc45;
// music[3599] = 256'hab433741c344884ff24f8a4a314b7a48d444ba4427432c4197436a4229348a2c;
// music[3600] = 256'hbb2f3b302830cc2c992bc32daf2b432a74287526f7232c20371b3a145c127410;
// music[3601] = 256'hfe0dd60e530cf5093a06d501abffe6fb6afa63f8aaf65ef666f371f182ef5fec;
// music[3602] = 256'h7be9c7e7c4e655e49fe260e026df16dec3db97d901d5d9d2e8d254d1f9d07ecf;
// music[3603] = 256'h2cced7ce5dcf1acc91c99fc9b1c6f0c641c74cc6dec80cc7bac795c81ec5bbc5;
// music[3604] = 256'h28c60ac61dc537c561c6a8c31bc5c6c6d6c644c663c5a9d16edd5edc35db56db;
// music[3605] = 256'h20dce8dc20dc99db91dc34df57dfc9dc3cde6be25ee1d7e14ce615e7aee828e9;
// music[3606] = 256'h6ce928eb37e9d8ec8beab7db8bd70dda19d9c7d9fcd90fdae7d962d99edbc7db;
// music[3607] = 256'h89db7adf69db48da6ce82fec5de97ceef9ec01eb36ed33eccbec82ed9becc1ec;
// music[3608] = 256'hfbeccceeaaf002f04aefecee82ee36efcdef24f16ff3cdf4dcf159eb3bece1f1;
// music[3609] = 256'hd7f20df504f6a1f30cf9930135ff30f952f85ef587f46ef7b4ed16e0d3e21eec;
// music[3610] = 256'hbff0ddf756ff0b023105d9070308c907c007fd076606ee043b04c102a0025703;
// music[3611] = 256'ha401f3017a0d3d187918971a421ccb1cf71ee01dd71fab2147239f2ad92f8e33;
// music[3612] = 256'hec37903a273c8f3e4042424492478549574bfa4d3b41b32b041fef1af71cdd1f;
// music[3613] = 256'h4222172481252827a7266e276b29e729a529c9289a29f82a652c1b2c9f298b29;
// music[3614] = 256'heb29742919291228ff27fd29f72cf42b2d290e29dc27f925be24b925cc29f929;
// music[3615] = 256'h8827f127cd260e24b22235235c285e2aa226f025a623af209620971ebf1e7a1f;
// music[3616] = 256'h951f37216320ad1f8f1f861f1120a81f4f1fcf1d941cb61b0d1a6f18bc15e613;
// music[3617] = 256'hd3102b0e4a0e410c2b099a063504b0ff3cff6d0a920f100bb008da053e03b400;
// music[3618] = 256'h94fdfdfbf6f934f800f69df483f4a3f2d4f0b6ef7ced91ecacec86ea9ee983e8;
// music[3619] = 256'ha8e5bde6ccdfbdd055cca9cccccb87cc6dcb99cabcc9a1c88bc849c773c6eec4;
// music[3620] = 256'h59c241c2abc291c142c087bed2bcc1bbd0baf0ba3abb4cba3bbac6bad8bad8ba;
// music[3621] = 256'h64bb64bd66beb0bd24bd1ebc6fbb3ebb20bb54bbdfb9e0b852baedbb1cbdeebd;
// music[3622] = 256'hfcbee9bfa0c008c2f0c22bc429c574c559c630c5c7c398c4f1c5b9c779c88bc9;
// music[3623] = 256'h66cbbecb8dccb2cd43ce24cf77cfb8d043d2d4d1c7d244d4dcd423d7e3d56bd9;
// music[3624] = 256'hbbe8d2efacee77f026f0e1ef54f0afefc2ef97f0a3f14af29ef4b7f666f869f6;
// music[3625] = 256'h2bef10ef97f3f2f668fc7ffe3afc77fed807e901e2eda1e813e83ce510e907e5;
// music[3626] = 256'h89d609d2fedb43e163e6faee40ef96f321f839f681f7e1f503f460f163ed19ed;
// music[3627] = 256'he2eba8eb60eb8aeafeeb0dee13f0c9ef52f2a5f5fff54ff8a6fad3fce9fe5501;
// music[3628] = 256'h9003bc042f081d0b3d0ee7104112b3144916c718e8190f1c941cbf1ea5338644;
// music[3629] = 256'h3f4429458a449344b4461f48754a6e4b214df94d604e804f764f86504e516652;
// music[3630] = 256'he7524a54bf546c533e5509534a57f966a26cce6dab6ef56a396a3c693967b466;
// music[3631] = 256'h9a66bb69b06cad6bc86a126af06641646663d668ea6d8a699269ba688a632065;
// music[3632] = 256'hdd5a8c4b114ba44b064c734dd74c834f0751e04fd04ee34ad646034618441d40;
// music[3633] = 256'h5b3d2a3b5639e135932fc1294d250f2239201f1eab1aba1711153911180f1a0d;
// music[3634] = 256'he60b620a98051d059afb08e34fd7aed6e3d39ed3c5d238d105d001ce4ecca3ca;
// music[3635] = 256'h1acae7c8bfc79ac63dc4e3c3b2c281c13ec2c6c091be2abea9be11beb2bde2bd;
// music[3636] = 256'h90bc6dbcacbba3bb0bbd21bcedbc7fbd57bd0dbe72bde2bd23bca5c19ed00fd5;
// music[3637] = 256'h07d329d304d344d3d5d28ed3b1d36ed325d4a7d40ed882d931d81ad857d7a6d6;
// music[3638] = 256'h39d7dad728d730d827d966d9d8db00d21bc5c0c619c731c645c8e5c736cb94cd;
// music[3639] = 256'h75ccbacc0acdf1cc55cc84cbc0caa2cb8ecc72cccacc5fcbebccd1ce66cc61cd;
// music[3640] = 256'h6ecd27cc62ce11cecccc13cdf9cd1dd1f1d298d2b8d3c9d3bcd1ccd239d41ed5;
// music[3641] = 256'hd7d8f5db30db8ed44fd1e4d600d9c8daabde47dd5adedfe5cde9a9e52ee1f7de;
// music[3642] = 256'ha3dbc4db16dbc1cf5ec653cd74d59bd9c5e37ae9a2ec4df146f007f10df153ee;
// music[3643] = 256'h51eb92e8cfe98ce74aeeb3fdeffea4fd57ff5d002d04e40480063d09270ab30b;
// music[3644] = 256'hc80e411287153d1c8d1e781cc61fe8212e24482774284a2cc93015349035ac36;
// music[3645] = 256'h56389b39253cb73db44066433544f7463e48a649454801472d4bee401f2f542c;
// music[3646] = 256'h932dac2c882d362e7a2f4c2f322dc72c0e2daa2c932b452bea2ec031ee302131;
// music[3647] = 256'ha22fa82b52295029052dcf2ff72d902dff2cea296728f526802bf03393314e2d;
// music[3648] = 256'hdd2b0d286d273a264d25a3268226e227ff279a273927f727022ace279529832b;
// music[3649] = 256'hb628bf28cd24af21cf1f751cff1d231bf3179f15e50f9f118f0e1c07d70b9c10;
// music[3650] = 256'h120e030a2703c6fb9ff8f8f305ef33f55afd67fc03f5cfe9c2e374e236de2ddd;
// music[3651] = 256'hd9e09de2cee1eee200e761e2e3d777d729d86ed626d77cd4e2d757db3bd80bda;
// music[3652] = 256'hacd4abce5ecfc6ceb3e068ef48e4b5df5ae207e263e4bde2bcdeffdb49db93df;
// music[3653] = 256'hefe3b6e35de319e433e130dcc8d586d239d9cddffde389e7dfe2a3dd2bd98fd6;
// music[3654] = 256'hd9e057e9c2eedef485e88edbaddae1d90fdb9bd1f0cc70d81bdbe2e6fbf8faf6;
// music[3655] = 256'h51edb9de92d582d8ffdad1e15ce8f8f1130218ff20f1edef7df4d0fc9b06ae0a;
// music[3656] = 256'hd20d740c7402bef961fb95fe25fac300400c59025ef7fe0130134a14d50ede12;
// music[3657] = 256'hb816111daa1c1d19f3294d33d22ec32a9d224a251522df1a9d29c82b8b1ef225;
// music[3658] = 256'ha32fd327e51f9027bc363c39a3353136452f4734c54167343923811b07126219;
// music[3659] = 256'h092dac3796313d22191e8c261529b5247d246a2823322b3424253522e4282720;
// music[3660] = 256'h0212ea1287262d3ae73ae12fac2e7329041f902bc22cae27f737d7359832642e;
// music[3661] = 256'hf220d8367e47a03ae02d33246e2cc92ccd1a981b4225ab29f12c7e249e0e39fc;
// music[3662] = 256'h2bfd53084f11e1143f0875fb67083c16e00de7f968e812e146e62bf7aefd04f9;
// music[3663] = 256'h63fc82f8f1ee74df4ad80af16bf840eaece32cdd6ce963f025df82db37e6f7ee;
// music[3664] = 256'h32ead5dfe2e4dfe8c8dab1cd4ed5fee28de5ecdb0ed1e6d6cadd73dbfcdf2fe5;
// music[3665] = 256'h6ee81beaa6de01d1c9d04eddedf295fc10e31ebebab7f0c96ccee9ca78d7cdea;
// music[3666] = 256'h3c00ddfaf0cdd5b46db98acc8cec3dfcf8092d1a4c0aa3e6f5cb81c83fd5d1e8;
// music[3667] = 256'he6f800ed16e248f64c0226f65af0df01101836212529a326da0e51021a051508;
// music[3668] = 256'h15159417fc053efb97f5eefefb22423bda39c539cd3a6c2de720f922b3242c20;
// music[3669] = 256'h8f192b12980c8b10d525983b004a7d540b48dd2da223602f2843b43f752c142d;
// music[3670] = 256'hb737873b49402b4bba5aaa5ede4b7538f035803a153e0a38c127f62875367330;
// music[3671] = 256'hca28802f3b332a24bb0335f174efdceed7f60ff450e748e444dbc5d4c2dc17d5;
// music[3672] = 256'hb4bcdcbbd4c827c514c72ccd39ccf6cb95bf32bbb9c8dacf3bd5c6d226c46dc0;
// music[3673] = 256'hd8ce62d6a2ca29c18eb968ba1bd09cdb78de3deb0df2d2e9e3d5bacd1ddd64f2;
// music[3674] = 256'h800344ff35f166f9cf0016f887f4a7fe790b03090606fe04bcf877f8f9fc4a01;
// music[3675] = 256'h300b0a041300f70075f98202940afd06890a1316d420081d4118121d811ec61e;
// music[3676] = 256'h711bc515dd1c492d95368c338327c7289839e936b031003adb3463361345b74e;
// music[3677] = 256'h19528b439c2f36267d256331fc3f7e49bd4c574a874c1655ae5bed5acc513348;
// music[3678] = 256'hd9438d40ca402640de34cc2a502f233aee355f329d3c353aa33b5b3ec22bbe2a;
// music[3679] = 256'hb637d939c83c413ea2364a211b14b5199a12b1045f0da71d5b18680979057508;
// music[3680] = 256'h1f0f6611ac0b94056d020e078a0e9f0ccd08390551f16ee10cebf6f3baf1c3e4;
// music[3681] = 256'h7ed987e40bf5c8fd04fd88fc6e04470020fc53fe7cf5d7f032f43aed4fe1d0e2;
// music[3682] = 256'he8e988e85fe21cd8b8d33ad5c5d7f1df4bdeffd012cbc5d560de24d09bccf9d8;
// music[3683] = 256'hced487cf3ecedec893cb23ce50ccaacbaec512c054bdf3b93cc339d336d791d3;
// music[3684] = 256'hd8caa8bfe0c173ca56c7ecc263be0caf4eac9abd56bca2a1a49c5ab0dab2a9b0;
// music[3685] = 256'hbeb607b76fb9f1b4d0a9f2a577abfcc023ce6ec8fac18db7d2ae70ae2bb7b3c6;
// music[3686] = 256'ha6cec3d2a0d161bf5eaee5b0d3b84ebfadc68cc64ccb22db4de4c1e696e1cbdb;
// music[3687] = 256'h2ddfe5d425c357cdf1e7cbf4f3f58cf8aaf6f7ef15f4adfbb9fd12ff10fddfff;
// music[3688] = 256'h2fff0cf155ea81f82c1add279e1eda2df82b1310180f4d179a1c3021a7247329;
// music[3689] = 256'h5e21a4211f316038bd34102fe52ee02c3830823e09458d446942bd3d3635c132;
// music[3690] = 256'h8c3db94264455b4b014c864ab6401639633f9042b541e14603515150c73e1839;
// music[3691] = 256'he744e94a404e06542452864a96446042b74491458c3fc23ad03a993c743e2e38;
// music[3692] = 256'h3c2ede2ba130a5399a357327922fd03e8933682a7f34682e7a2a9b35b52b3a29;
// music[3693] = 256'hda2df61e881f73239322522461182c19331d31141b11c50cdf10fc13e00a0d08;
// music[3694] = 256'ha7068e0fea1c6e19d51382108d0fec125213420ec8094c0e240961fc88ffeeff;
// music[3695] = 256'h5efa0af518f20e0197042e02b811ce09b900ff0ba5099511371ac30e390c9406;
// music[3696] = 256'h5203830cd6087809df10ee097404110281fd79fe8900cbffd9f90cf7e5f841f3;
// music[3697] = 256'h64f9920223fbaef9e0eae0cd32cd75d94fdba0d64ed7e3da18d11ec9bbcfb6d8;
// music[3698] = 256'h35d790d149cf44ccabd640daf2ca4dcb73ce8ad35add15d3f4c9f5cd5dd216ce;
// music[3699] = 256'h0fc584cb0dd7eaddaed990cc30cf5dd6aad679d70ed30ccfebd29bd75cd65dda;
// music[3700] = 256'h37e257dd7fd666dbede246df50da8bdee5dd42dbfadd25e698eadcdea5dd6ae4;
// music[3701] = 256'h6eda1ed5e3d975de03dfecd59ece2ad231dee0e61beae8ed3ae82be2f1e684e9;
// music[3702] = 256'h59ec15f2a1f383f322f33df319f4e3f235f302f62ef5fbf031f3fffe1704a4fa;
// music[3703] = 256'h06f3eaf54500470799fe21f836ffc1004cfec9fd5501600f8a103903c1ff52fd;
// music[3704] = 256'hf5f5bdf3f001860f0107ee034b062008b8164e12b6055b08b00251fd65016704;
// music[3705] = 256'h7f07ed087800a2f94a06a20bfe05b6086f062407b00abe045102a3036004d804;
// music[3706] = 256'hc40563087f09a5ff45f8020cf414910a5b0ff80ec60dea0f24068f09b0120e1a;
// music[3707] = 256'hac2b03306e26c32678290328672cc530e62c6f2595238d29342e453474301526;
// music[3708] = 256'h382c482f802948296b332f400137432d562ac2257b2e24331835eb36f5301231;
// music[3709] = 256'hdd2b5025b423d425c22cf029cd2aa72bdc25c22a092c382b482bce239f205c23;
// music[3710] = 256'h342b8d277a0e0b000606dc0b990d790e900bba076c07650895075006cf070307;
// music[3711] = 256'h5e03dbff0afffb07f00c7f078e08040a97084c0c9d06a1f9bdfcfb07b60b120e;
// music[3712] = 256'h6910550bf6020603dd05b803b604bd076f04d3fead062810c00c62133e16b40a;
// music[3713] = 256'h9d0bfa087202d806bc0c1814d110e00a1b119c0cac055e0cd70b1105ef06d90b;
// music[3714] = 256'he313b21440087005dd0850091b0ff20e02092a07db0496026a048f0a6f16571c;
// music[3715] = 256'he7103c063b06bf053a04e1070e110b0e6607030bdf0419024d08d0068408ab08;
// music[3716] = 256'h2f06e207f50a7d0ce405c600f7ff07001404af04b9048904b100d7ff9c008502;
// music[3717] = 256'ha70a900bde008d09b91b9a1eb12196201c1d611cc6180f1bb414fb0b6a10c419;
// music[3718] = 256'h191f9213c00d2a1398105e10670972050d0f1b103e08b603b30f8c19700ac0fe;
// music[3719] = 256'h9a01300679075402cdfff306550aa20673049ffe88fcc7fff500110b6c0d5009;
// music[3720] = 256'h9111e612b210670e8e0b0b17e0179806d30035064b04aefd240084002cfd9003;
// music[3721] = 256'ha607b7071b0701feedf67bf6d0f75cfdd0000afb04f3d5f077f1abf4acf512ed;
// music[3722] = 256'h61ec41f274eb54e7bcee18f473ec86e186e6eae602d8b8d231d640d820d6cdcb;
// music[3723] = 256'h16bb7dadbab0b9ba01b409a7acab90b154ad45b2a6b15ea89ba917a769a7d6aa;
// music[3724] = 256'hb0a4d2a6a2a968a67fa681a6d7a9eaaaa7adb1b1dfa74f9e019e8aa2aca8d3a8;
// music[3725] = 256'h0aa5e8a536b161b5dfac08a836a12ea2adadbfb3a7b76fb382aaf4a7ffa528a5;
// music[3726] = 256'hf2acf3b8d7b3edae20b726b3c4b0c4ae96a947b114ab18a470aebcb1edb100ad;
// music[3727] = 256'h22a6fea72faa3eaee5b0d0b22bb45aac48a739aa80af68b252afb5b332c08ec2;
// music[3728] = 256'h78bf26c09ebc6db5c0b41fbb6fc17bc56bc8f5c607c3f8bf30c214c8f3c5ddc7;
// music[3729] = 256'h52d133d207d39ed1f3cd5fd2d2d2ffd315da2fd8ffd310d816e201e268dce4e2;
// music[3730] = 256'h27e6c0de77ddfae691f135f39cefefeb8ce8d5e8eceb52f2abf659f226f280f5;
// music[3731] = 256'h05f263f3e3f643f51ef8edfa07ff3106d60579069306b90058048c0ec012450f;
// music[3732] = 256'h29079505fd0b280f961041141a0ffb0df71eea2111182e25a7365e36c636463a;
// music[3733] = 256'h72363338513fef3b80378f39ae397736443cf4473543ef42654edf45df3f5747;
// music[3734] = 256'ha4494349d0411d44e94f7f4d024a3b469143104cfe53bc5658502f4b70519d54;
// music[3735] = 256'h9156f9534b49cc46be4dc3584a5b6256ce5a4a59054f964a3b4ef0580451f33c;
// music[3736] = 256'h313dd03f823bbc3a4c40904c5d4f2c4a124b854d664a0e45fd47c94ce94be049;
// music[3737] = 256'h8f48de486948a54882481745d93f784324540552c849e3528e4dbe4a224f7648;
// music[3738] = 256'h5c4d0e50b551d0573f4bae44c347bc47c84d5a4c384af04ff54a564b5d56f552;
// music[3739] = 256'h4952ba5e2c621f6152608b5f91610b5d7d51c74c18513f51a4507b5203513b53;
// music[3740] = 256'hb750944b864adf4ca950fb45cc48d3569a4f3b54ce57c44f454f8f434c42314a;
// music[3741] = 256'h9f46f94859468b3f68418941c83b9e384738c23240379140413c4b3432308e38;
// music[3742] = 256'hf73c2a309d306f3aab39a135dc36c23625307f30e62d3d243027ca247621b72f;
// music[3743] = 256'h6730d225332602222e1faf228f1a8813d619221d3f180715a2147f12bf0dc003;
// music[3744] = 256'h7000c709940b00055dfe97f9dff944f3a7e77de28de3fce8f9e9bae393e015e9;
// music[3745] = 256'h8ceedbe26bdcccdfa9da2dd5d6d858dd59e409f10bf445f250f3dfecebec95f0;
// music[3746] = 256'hfdeb94ee2ef095e877e547e893e43bdc85dea3e032da48d773d6f5d63ed880d7;
// music[3747] = 256'hcbd6f4d3c1d110d638d772cd6bc7f0c92bcb86ca12c624c758cf5ccc03c430c2;
// music[3748] = 256'h83c382c335c0d2bea3bf18c2d0c48ec0d8b841b4bfb700bb83ab069cb79d9aa1;
// music[3749] = 256'he6a2549a8693df9e75a0ce9b049c1295e19a059fb695b89ab79d94990798e393;
// music[3750] = 256'he898cb9bd5947993819513979496ed9320948e966b978a98059bd4980d972196;
// music[3751] = 256'h1797939ee89b65976b9d5b9ed39dca9de49d5fa0d0a01ca1be9d249e5ca769ae;
// music[3752] = 256'h84adb3a35aa217abc8adefaa7ba474a1f7a203a82cadafa96ca6d5a79eac1cae;
// music[3753] = 256'hbfb00eb983add5a82ab3e2abbdaf15b6afb1e8b66db312b7cfbe9eb331b59fbe;
// music[3754] = 256'hf7bb17bd66bd56b84dbb03c1c9bf42bd6abc0ec379cbfbc953c7d6c7b6c92bca;
// music[3755] = 256'hf4c678c919cda9c8cac61fcbaaccc9cc18cb0dd058da49cedcc661d249d07dd2;
// music[3756] = 256'hfcd4d2d139d938d5bbd1a7d618d633d584d151d30ed8e3da59dc71d587d260d3;
// music[3757] = 256'h4fd51ed67fd781de82dc50dfa8e913e8b3e742e630e135e73ef2aeee0ced69f6;
// music[3758] = 256'h2ef195f01bf547ee68f19ef27fffdf175a193b192a1b0d1941194b16d719fd1b;
// music[3759] = 256'h6d18b019d51d0f200221c524f72443221d20b923ec307730142a2c35053cc734;
// music[3760] = 256'h9030a82f5b32a63df640003b64363d39e14ca65a615b0859dc53055fcd614254;
// music[3761] = 256'he45b32659d60915fe561be621860395eb75f1157f646be4c9f4f9e42ef4cad4f;
// music[3762] = 256'h9441e746cc473944814b8b503d4eef495049e94629449144414700520b586750;
// music[3763] = 256'h94473e458947eb4f7555c851b7518951194fcf51465168502e53c5555652014c;
// music[3764] = 256'he44b254ea057f260605de6597a54314da352f55d4d5d2e580b59fa58cf5c8f5a;
// music[3765] = 256'h494d594fc75d9661cd59135cce5dc451d7559f599953c952204c1453c3569845;
// music[3766] = 256'ha0415341903fad40fe3ab3371d395e3c5e3cda3c59454c45fd3b9f37ce380b3d;
// music[3767] = 256'he243df464f3ede34f936833ae6387239214069493d494b3d09368538a73e683b;
// music[3768] = 256'h7330d0392e4ab5433d3cb23fa43b733657398238bf3aee3df439f03ddb3a1e30;
// music[3769] = 256'h8134493783374c383a321a2dfd29652d9a30242e52313330f52bd72c21264b22;
// music[3770] = 256'h1e2d4a2e62254022b91e112122240f1ec41daf219f243a1fe211a2131f1d111b;
// music[3771] = 256'h4015e718561aac16a023f92d332a61285d23982472279c25c227991dd614ec1b;
// music[3772] = 256'h931b65176f19431b6b1b3b18c00ff80a0b0fca10470e3c0b8f09190be7036401;
// music[3773] = 256'h9e0d970a8902b7038ffe25ffff0397013cfe5ffdfa009afdc6f6b5f8fcfbadff;
// music[3774] = 256'hd80279009cf4ffef3ef8f6f574f67af1abda7cd73eddc7db3fd91ed2c7cf44ce;
// music[3775] = 256'hbecb68cf9dd4e1d289d02cd877d308cc67d078cedbcc13c808c73ecd3ec761c8;
// music[3776] = 256'h40ca72c15abe95beb6c131c037bdabc207c3b2c10dc378bd30b810bdefbe01be;
// music[3777] = 256'h23c5bcc259bb63bffabfdfbacfbba0c09cbdd3b6d1b872bb36b8d9b713bb7ab9;
// music[3778] = 256'h37bad4bd59ba67ba1fb966b086ae5caf69b008b2c4aeaeacbbb004b2a4adc8ac;
// music[3779] = 256'h28aaffa875ae6aabbfaa15af24ab7fa914adc8ae6dac6caac7ac25af4eae58a9;
// music[3780] = 256'haba958ab3ca780a8f5ab5eac7aaca3ab36ac92ac5fa931a4a4a588a98faaccab;
// music[3781] = 256'h4fa6d9a2b4a589a36b9e9a9a9ba1a9a7bba20da437a13c9ba2a105a567a1459f;
// music[3782] = 256'hdd9c6d99d59f27aff3b3b6b483b5f3ad03aed1b5ceb558b1b8b07db419b341af;
// music[3783] = 256'h94afdaaab3a967b37ab6b6b39cb240aeccac9faf11ad93a9eaaae6ab19af38b3;
// music[3784] = 256'hafac53ac79c185cd54c8f6c9b0cb8fcbe1d2afcf4fc674cb0bcdd0c45ec931d2;
// music[3785] = 256'h90cfc2cfa4d539d35dcd21cf82d388d215d2cfd8d2dc33d8e3d40bd5fad58fdb;
// music[3786] = 256'hd7e07ce058e070e34fe7abe593e1ede13ce027e297e851e5e5e553eea4ebf7e5;
// music[3787] = 256'hb9e714ea0ded30f00fed4be33fd5c5cba2cdd0c82cba8ab803c2f0c6a7c23fbe;
// music[3788] = 256'h32c2ecbf84b6edb8cfbf10bdfebb24c4f8c766c551c3c2c204c6b5c43dbfd9c0;
// music[3789] = 256'h1fc572cbadcebdcba1d03cd218c73cc597ce97d248d35bd467d2e5d31ed72ad5;
// music[3790] = 256'h05d522d578d401d9fcdb99d816d7ffdafddbdfdba7dfc7dffedbd5d829df8ee6;
// music[3791] = 256'h82e13ae436e927e581e720e529e42eee6def6cec6beb27e711e635ec60f06cee;
// music[3792] = 256'heaf10ff547ef89ee74f547fa76fbeefc6afeadfe42ff20fff1fd10ff26036c03;
// music[3793] = 256'ha003140a610a38063707e60c9c11880cd809c10e7d106512ac13dc161d1b0618;
// music[3794] = 256'h7613e6118b13581692161e18d31d9421d31cd21bf622e524e621ec1d4c1d9b21;
// music[3795] = 256'h8d22f322d925a8262528d5298d2596252e2ffe2fe329c92bae2e7e2be5263227;
// music[3796] = 256'h222acd2bc42e9e2f0b3008354d34be2cc72be332d8374a34b234d93ceb39583c;
// music[3797] = 256'hff50905707549f58dd598a5797563b59d65ce7596d54675343584f5915562459;
// music[3798] = 256'h075d5e5dc45a575a31607f5dc157f75a465958589c611c65a0615360625ba256;
// music[3799] = 256'h785dc86429634d5f035c035cd15c4e5e5c63ad61505f9c63b3624e5d2f580a59;
// music[3800] = 256'h625f3e61905d794fca42e444c044144042426a48bf46883eeb3c283c633b453c;
// music[3801] = 256'h3839c739cc38ae36423b8f393638223d5e38233190321e3248302a36493a2035;
// music[3802] = 256'h403175333d351633772f652c812a282c003383361d330f35a137b33327320a2f;
// music[3803] = 256'he82e0935c333bc30db2cef279c2db0319b2e7a2d4f2e4331e43297381c426a44;
// music[3804] = 256'ha3450e439d3f9147ff4913438b41ce43b240d939483e3e43303e693d2c3de63c;
// music[3805] = 256'hfd3d7b3b753c183d443eac40c63fb641503df835cf3b3a430f40163aaf3ca63d;
// music[3806] = 256'h8f37e839fe3deb3d6a3e123a19381b3bdd3899379b3c743ba432a72fa531f131;
// music[3807] = 256'h792faf2cb52e91309c326e34f42d482b242b46247825a32b922b5b276a265c2b;
// music[3808] = 256'hdb248b18131cdd250627ae22e1240426c6204921d11fd51c631b3e1607172a17;
// music[3809] = 256'h3c148317da1a5c14b00010f593f715f8f2f6ddf25cf010f0d9f0fdfc67047305;
// music[3810] = 256'h390dc20d5109fb08ec0761073406af051c04e4fe0b0075010cfa67f7d6fbeefd;
// music[3811] = 256'he1fbf4fb54fdf2f699f207f348f197f3c7f2aeeeaced03eee4f28bf279ed4fec;
// music[3812] = 256'h12ea43ecd3ed84e839e88ceaabe8b6e88de9ade59ae249e02bdd44e091e3e5e2;
// music[3813] = 256'h0edd49cc19c06cc12fc108bcd6b966baf9b74db34db457bab3bb82b944b950b7;
// music[3814] = 256'h1db524b55bb469b211b0d2b2d0b7b5b35eadddac32aeb7ae91adfcaed1afacac;
// music[3815] = 256'h6aaf12b179ab4fab4aad99ab6eac7eaed8ac1dab5ea9f7a671ad5bb120aabda9;
// music[3816] = 256'h22ab0babd9b05eb293ae3aa897a31da602adc5b138ab20a6c2a96eaaeeababaa;
// music[3817] = 256'h2baa1eb0d5a8c79d87a32fa8d7a720af2fae03a6b1abbbafcaabbead66ade6a7;
// music[3818] = 256'hd2a50da742a8a7ab0db150afc1ab11af53b2d0b1beb09ab0d0ae96ab77ab31ae;
// music[3819] = 256'h99b10fb267adc5abb0b189b3ddaf28b02cb045b069b1ffad62ad9dade5a9d7aa;
// music[3820] = 256'h51afa4b27eb268aeddaadaa85daa1aaf5faf52a9b7a715ae83ad75a826ad8db2;
// music[3821] = 256'h2ab234afb2aa53aa1dab08a87ba7d0aedbb474aef8a8faaa02abc9ab91a905a7;
// music[3822] = 256'h81aabdaa3dab7eac2aacfeadc4ab4cac12b16dad7fac0cbb4aca53ce65cfc9ce;
// music[3823] = 256'h05ce97cf75cc59cdbdd06ece81ce58cfa6d18dd391d177d160d05cd191d223d0;
// music[3824] = 256'he9cc4dcff6dd07de31d3bcd751d6c1d75adf6cdc80e08fdf62dd3ae370db20dd;
// music[3825] = 256'h1ae4eddcdfde2ddf8adee9e5a8e058e41ffada0099fe6700c3fd3efee3fd07ef;
// music[3826] = 256'h07e7e9ed0bee1eea71e89ee610ec29f013ebe4ecc5f233ee37ebcaf4c7fd60fb;
// music[3827] = 256'h8ff833f79bf1b3f64afb8bf60dfccdfa4ff690ff2901e0020f05e3fd02fe2bff;
// music[3828] = 256'hd0fd5bfe0afe4702df0575073a073a07740ed60e37075e08ce0cf00a880a9911;
// music[3829] = 256'hf812e10e751423165c0c650d4f17bb158b10e917801d8e173818551b33193f1d;
// music[3830] = 256'h551e4b1d4d1f2e1b891cea204520c123542454227021101e7920f825ff1f3012;
// music[3831] = 256'hfb0e0f125b10cc13241758147217031dbc1a6615fe16031c351f7b209b1bff1a;
// music[3832] = 256'h44248f268a23262482220f24162ab826ad215223bb24ed289c2ab728ae2d5b30;
// music[3833] = 256'hc92ddd2af0269d251027a72f87338a2c9330bb31812c2433f433a536463b4a32;
// music[3834] = 256'h8e34473a97370e3aba37e032b832a235d4372e336030af31883684392f35c034;
// music[3835] = 256'he233f931fc33ce32b434f2372d38cd3766379942d150bc4e9a4e335866557d50;
// music[3836] = 256'hd055e854425374536a51df546f5525544154dc4e4f4dfe4f6251ca524a51374d;
// music[3837] = 256'h64494048c84ab44ad447ef4bc34fb44ce54eb550004e764d254b164c1a4fa44a;
// music[3838] = 256'h59476a4bba4df44a9646944274430345ab47004b374347426943df31072c2931;
// music[3839] = 256'h392c2f289024132210237123f3228221d71e4b1d5a22ec24d3223f25d821321b;
// music[3840] = 256'h891b0c1f762271238021741d421ec121821e491d161c5518261c331eb5187616;
// music[3841] = 256'h981853195217a7171a1d3b1f741a97180b1a9919111808144a12b017601b0b19;
// music[3842] = 256'hc8180d1b9c195a1706169516931920172d129111a4112b1271147116be154f15;
// music[3843] = 256'h2b194319d9115911ac19b0182614ff17b21564104a137a1461148516f8163716;
// music[3844] = 256'hab14b7139f14fc156614c610e0129c178516be13b815c719561a571730137412;
// music[3845] = 256'h34181918e50ed40ee615c016e9145c125211e712c8123e134b112c0e230f030e;
// music[3846] = 256'hc30e9612cf127d124d0f9c0ab009a70a970b560ac10bd00d3f0a0f097e0ac10a;
// music[3847] = 256'had08d608e9166021661c311b971a9c1a9d22931f1f177a1af41c6a1974146913;
// music[3848] = 256'h1118c717ce12bf10fd124314c5146b21732da02be729812719247127202a0c28;
// music[3849] = 256'heb261c27bb249425b0269c1ff01c7b21b223b823e120e01c0b1b8b19c6178b1a;
// music[3850] = 256'hc61dfe1ba11db51e3b1d291cb114d912d4168b16b01806175113071213115714;
// music[3851] = 256'h721308138b146510351344151411df0f500d300c510357f3c5f0f2f17ff16bf4;
// music[3852] = 256'h18f41ff547f42aef97f00ff07fec42f093e93cd753d21ad8aad7a7d1b3d2bad5;
// music[3853] = 256'h44d151d385d5f6cfe4cfbdd00bd29ad34bcfaecd1cce03cef3cd0acdd0cce5cb;
// music[3854] = 256'h57ce72d3f0d4e1d1bbcfbcd10cd001cdc0ca77c7f5c810cb1fcc2ccc4fcb09cb;
// music[3855] = 256'hf5c7dcc514c862cf3dcfb2c8e4d063d3e1ce88d086ca14cc9cce3fc825cc22cd;
// music[3856] = 256'h89cdc0d254ceeac96dc914c766c65bc845cb11cd0cce40ce77cd4fcd09cffcce;
// music[3857] = 256'h49ccf5cb4dcd68cea8d14fd672d75ed61cd718d792d728d753d501d66cd8cedc;
// music[3858] = 256'hfddc1adb59dbf1d692d8d3dd4fddbedff2dcd2d434d4c3d86ade6adeb3d818d9;
// music[3859] = 256'h00dc24dae5dbbddde7dbbadf94e03edd1fde55df0fe2cae236df9fdce8dbd2dc;
// music[3860] = 256'h9cdc34de7edf75df9be215e166dde1de7bdefdd925d931dcfcd9dfd80ada93d9;
// music[3861] = 256'h40dcc7d931d6b2d878e065f003f866f88bf8a7f043ed2df097f1fef38ff6c8f5;
// music[3862] = 256'hf4f06af143f321f264f588f536f285ef17eee8f014f1beed11ed14f1c7f441f2;
// music[3863] = 256'h66ed6beca1f130efb0e93ff1b2f3e5f1dbf1d6eae1eb03ee4ceba6ee66eefdec;
// music[3864] = 256'h50edc5ed4def97edc9efc7ee03eb32ed3be05acd4bcd95d553d75ed201d32bd4;
// music[3865] = 256'hf5d0e3d3ccd3ffd233d5b3d0d4d032d3add034d2e6d1c0cfd4d0fecf89d2e3d7;
// music[3866] = 256'hddd5aad123d1b9d4aad9afd478d0ccd5e6d42dd20dd381d046cd7ccc77d0fbd0;
// music[3867] = 256'hefd000da16da9dd1d3d16bd4b2d424d495d1dace81cfecd160d2e0d27dd272cf;
// music[3868] = 256'h18d11bd826d907d649d6ebd6b9dae4d95fd26ed8a2dc48d60de07debdbe9edeb;
// music[3869] = 256'h8ced41ea90e915ec57ee89ea03e85aed04f097ef9af0aceeb1ea12eae8ebb0eb;
// music[3870] = 256'hffebcaebcfe8cde9daebede9aae8a2eb5def80edc9eb22ed46ec3bec95edabed;
// music[3871] = 256'h96ec1ceb26e938eaa0ee66eefaedb0ed9cecadf047edceea7cee05e942ea8bef;
// music[3872] = 256'h3cec26ededee4aeeb3ed50ee2fefe0edf8f1b6f3f2ed73ec04edfeee5df2aff3;
// music[3873] = 256'h93f36cef96ee66f301f419f46df482f39cf4fef019ed9fefb3f1c7f17cf019f3;
// music[3874] = 256'h4bf206edd4f80a00c7f7fdfae6fb75f745f9d8f84bfa61fa99f828fc37fd32fe;
// music[3875] = 256'h9b01a5ff68fc02fcd5fb91ff0702d5fcf7fbccfeae00b403520175014b057603;
// music[3876] = 256'h5704a9054104a404aa02d5018f052908fa0640051606d6066008760aa90a340c;
// music[3877] = 256'h820da00db50b1808a70c880ee5ffa4f3f8f3fef637f7bbf255f2cafa88fb73f7;
// music[3878] = 256'h06fe410005fe6d00c4fa21faa100edfe3d01920217ffb30025036d05750196fc;
// music[3879] = 256'h7b01df037f028703960341018201db04be04d2037a05520765068f03f306040b;
// music[3880] = 256'h220afe080b0788076d0a0709ec060609ca0c310f490f2610421340117f0e540f;
// music[3881] = 256'hbc0e6b10740ec20b4512e313a012e6141e13501162129813b811c211c9178218;
// music[3882] = 256'h61157715c515f1168118c0187019b41a231baf1aa418bb16c218a11d0f237124;
// music[3883] = 256'hce206c1efe1c781de022c126f92558273f2ab928ec27e42868263e2546270228;
// music[3884] = 256'h3528c42aee2a2328702873285c290e2ba627e927eb2a102bff2dee2f6a2d482a;
// music[3885] = 256'hb929af2be92d9f2f8f2d6c2c912e9d2c122a09294b29f82c102d8a2b902c3a2c;
// music[3886] = 256'h6d2c7a2da02f3930692c262d3e30f02e252dc92b272de82cab28502b4b2dd629;
// music[3887] = 256'h013346413a43e345114b3149b8489249bc467f438644a34992499e4b9a4ecf48;
// music[3888] = 256'hca485749ca478b4d174cf949674c9b498149c349b547e148f948d948f0495447;
// music[3889] = 256'h7b456648b4484a488848d74547449644f846ea46914515488f469145c746c547;
// music[3890] = 256'h234b2149c248bb44733274272030c53feb44d243e843b941d9441a45b5426a44;
// music[3891] = 256'haf418d429143c43f70408342b445ca459b430c420f3ff5404c420340ff40bc42;
// music[3892] = 256'h5641433d763d2f40f53fb93e723d253d793b233b633e243dab381038db391a39;
// music[3893] = 256'h9237a73708397639cd365e39903a503545387639ed355637a834ab3280323530;
// music[3894] = 256'hdb33d43669339931cb322433b332f731f9304631a630c430f330c32d842cbf2d;
// music[3895] = 256'hcd2f6c31672eb82b212c1f2b5029962cc72fa12c4a2d9e2f352c9f25d719f713;
// music[3896] = 256'ha316351547162b193d16f21381138e16801aa915af10aa121214ef136712f70f;
// music[3897] = 256'he30e010d6c0bdb0cf20f0e107e0ddd0cde0b050a7909fd09f60a1d0a5909f008;
// music[3898] = 256'haa07bb055b05ee08d405d900a804040249fd24005f019402a20140fd7dfc43fc;
// music[3899] = 256'h42fa45fa4ffd49fcbbf7d2f85ef80cf31af5dcf8f9f6ccf672f188eb57f9250a;
// music[3900] = 256'h410d7e0c020b040b9b09d4052506110652059605f10526072705f6022203ef04;
// music[3901] = 256'h4d0644022700f8003d00f400b6fdf7fa23fd5cfbcbf9aefa42fa57fc79fcaaf7;
// music[3902] = 256'h86f6f9f845f94ef9acf7d6f3bff205f3d9f37df37cf239f38cefc1ef18f312ed;
// music[3903] = 256'hdaeee6ef34dee5d246d222d287d40cd45cd25dd084ce3ccf02ce72cdabcd3ccd;
// music[3904] = 256'hedceccce5bcd4bcc33c9a4c827cb4acb30cb65cc3ecb5ec900c9e0c9cbcab6c9;
// music[3905] = 256'hcfc765c7b0c9c3cbafcad7c7f0c3e7c309c60fc52ac527c5ddc249c040c05cc4;
// music[3906] = 256'hbfc4e8c118c26cc26fc109c20ec380c054c05dc185bd01bf71c25cc19ec0b3bd;
// music[3907] = 256'hafbcbfbdfcbcbebe24c2e0c3e1c0f2bdb5bf3ac086bf86bd35bba9bb2fbdeebf;
// music[3908] = 256'hf0c082c00dc266c18abd75bc7ac180c325c098c007c149bf34bf29be7bbd7dbe;
// music[3909] = 256'h6abf4cc14ec5e7c523c1e7c00cc447c6cac842c6dfc471c60ac35fc147c205c3;
// music[3910] = 256'hb2c32ec348c61fc61bc2dcc3d0c32ac1e6c1d1c178c068c336c873c448bf51c0;
// music[3911] = 256'hf4c08dc374c2a6bc88bf27c480c4e6c31cc355c5a2c480c1c1c1eec0b9c2afc4;
// music[3912] = 256'h5bc23cca4cd6bdd613d59bd4c3d327d547d675da02da04d7b2e580f3cdefb7ef;
// music[3913] = 256'hd8f7fdfc3efb0ff85ff862f6ecf407f76bf5ebf445f9f2fbd9fd190034018002;
// music[3914] = 256'h53027b01d90274044a037e02e0062e089903dd0316058303e903d702a6002800;
// music[3915] = 256'h4f00310062ffe7fefbfbdbf92dfd96fd0cfb49f9c6f433f31ff42cf41af8fcf2;
// music[3916] = 256'hd3e2bedd2fdf58dcf1db78db16da6eda7bd8c5d6d9d823db69d98fd78ed954d8;
// music[3917] = 256'h58d6bdd824d830d904dc92d9e6da33d865cafcc4c7c67fc51fc733ca45c9bdc7;
// music[3918] = 256'h22c964c9c6c70fc8fdc858cbc8cc2acbf0cb36ce76cf20cfbdcc11cde7cf74d0;
// music[3919] = 256'he5ce00ce1ccf8bd1eed26ad1c0d219d865d739d4aed5c4d4e0d4e9d905da50d8;
// music[3920] = 256'h5ed97bd84edbcee04cdf7bdb71dc9adedfddb2de65e2bce22de3d6e66ae7a8e6;
// music[3921] = 256'h0fe7b2e58fe5efe6fce7b7eadbeb50eb8cec58ec45eb51ed2df23cf63af8c1f9;
// music[3922] = 256'h61f8bdf64df8d9f842fbcafe64fd19fdc8ff8aff9cff3a014300adff2900b4ff;
// music[3923] = 256'h07017302fe024d0484045b023a027b070909f7069d096b08a606b80b170b2007;
// music[3924] = 256'h9008a907740571064b05aa04f2067008c10a860a7d08410a4e0ca60cdf0bce0c;
// music[3925] = 256'h7a0c9e08470b420fd50e540e780ca30dd70db70fa41d7a264d248025c127d327;
// music[3926] = 256'h9c284e284529bd2c0b2d1b2e7230d32d6b2d22302f30dd30fc31dc30982ef430;
// music[3927] = 256'h4934583123315a32602e0e2ea52f1e2f9830cc31c531c130882fd83040311831;
// music[3928] = 256'h403281312131a3313330342eb92e7c3257333032a9339834b334af2b231cc31a;
// music[3929] = 256'h701d6f19a91a101cca1bff1d401c861964182e1a511e8e1cb11c4f20c11e2b1f;
// music[3930] = 256'h7a1f691eed20da1f471d3b1d7a1d4820fe221c229b20ce20861f1c1f2e20241d;
// music[3931] = 256'h401c801ee21f411f31189d169f1ba41a1f1cbd215a233122ca218d21501f091e;
// music[3932] = 256'ha01c3e1a7519291708160418111819167e159415d9143b16a018a7184a19991a;
// music[3933] = 256'hb81a481ad019761bb31f5d223524a5251925c2250c242d27bb36323d653ba63e;
// music[3934] = 256'h3940c042c0432f42d54443462f48bb4aca494a4a604ca34c3a4cde4cc34bed49;
// music[3935] = 256'hc74aa94b6a4cd74c8e4d754e4a4c514b424c6c4b2b4aa948844794461e449642;
// music[3936] = 256'h76433c435841c93f793faa40e33e553cd13d9f3c07389c3676377d365834a932;
// music[3937] = 256'hc92f112eaa2d2b2c262c082eff2dae2aa5286a28902838294f25be2298237b21;
// music[3938] = 256'ha820a02068204b1fd41dbc1f631d3020732e43351d34ac322f30f92fe431ab30;
// music[3939] = 256'h782e512f5b28731bc71681163d16681570140b152b1306116010210fba0e860e;
// music[3940] = 256'h8d0d5c0b810a190cbf0b280aac09b7092809a006da041906bd074a0777067a07;
// music[3941] = 256'h9f060d04e00302036503f604b6028002ac01660020025cf60de738e7f6e987ea;
// music[3942] = 256'hcfe964e702e8c5e731e6efe4cee400e65ee4f6e350e612e533e34ce48ce4bee3;
// music[3943] = 256'h1de48ee360e24ce22de3cee3f1e208e394e3f3e235e348e493e5ace44de3aee3;
// music[3944] = 256'hede14fe11de3ede2e6e2d4e325e3b7e1e1e27fe39be1a2e273e3bce1c3e195e2;
// music[3945] = 256'hcfe27ee23ee3b0e456e4fce35ce40ee622e732e56ee49ce405e5f3e695e6cce4;
// music[3946] = 256'h8ce4d4e55ae872e947e825e814ea85ea84eaefebf8ebf8ec64ed58eb90ec72ed;
// music[3947] = 256'h9feb3deb7bed9aefceec71ecabefb6ee2bf0c1f19aefb8ef49ef53effef08af0;
// music[3948] = 256'h41f0bdf056f1dbf174f177f1c0f37bf62af562f253f207f325f398f396f362f2;
// music[3949] = 256'h07f242f1f7efacf0a3ee51eb88eb20ec31edb5ed05ed7eed0cec52ea8aeb22ec;
// music[3950] = 256'hceeba3ec02ede6ec2feda1eb77ebb6ef95efceeafaea29ed4ded87eebaeebded;
// music[3951] = 256'he6ed9bec3fedfaeeffeb28f2a20212087f06a6068803540375063c067a046b04;
// music[3952] = 256'h5c0700086106c9076f074506f30603061106c9061b06e0068d070e066f050306;
// music[3953] = 256'heb048903d903e1055106ee036e0479051104cf0322035e04c206dd046d036a04;
// music[3954] = 256'h1a03510281056705c9038205d803c104cd03eef498eaeeeb2eed4ced2aee0bee;
// music[3955] = 256'h2cec86ecc0ec00ec9bebdbeaa1f5b9010401e101a103e801e501a00174026c03;
// music[3956] = 256'he2023e02cb012e018f0066006fffcffe03000e03500422038f049d02b900c203;
// music[3957] = 256'ha402c302ea02cf000403ad01fbff75012d00cdffb8ff4600fe00a4ff76ffb4ff;
// music[3958] = 256'hf6ffc4fff9fd31fd24fe46ff4fffd7ffedff41fe4efdc4fd4ffffb008a023c03;
// music[3959] = 256'he7015b01a3002fff2801e603b801baff4601cdfffafea201040148006600f9fe;
// music[3960] = 256'hc5feb9ff780171024f010001a802af023c0123029e026b028afd00f1a5ececee;
// music[3961] = 256'hf5ec22ee04ef4bed80ef51f172f184f198f01ef021ef5dee1fefbaeef2ed43ed;
// music[3962] = 256'h75eb2eeaf1e9e3ea12eb55ea48eb9cea56e923e9d1e7a8e7f4e770e81ce8dae5;
// music[3963] = 256'h1de7bae875e79ce765e88de704e7cbe7cce660e6a3e94eebb9ea30eb33ec70eb;
// music[3964] = 256'h5eeb28eb68e9b8f3b20246036302ae044e024c00b8ff1c00a00186029102f601;
// music[3965] = 256'hfe01dc010a024b02b0018403c50564050404690210022e02cb0093ff60007801;
// music[3966] = 256'h6a0044009a01840061ff3bffaafe89ff56006cff2dfed9fdd5fe2a00de00d400;
// music[3967] = 256'hf300caff38ffcbff85fd19ff03fde7eca4e4d7e64de582e59be61de6dde588e5;
// music[3968] = 256'hb8e6e4e6b5e573e5d8e6fbe7cce647e643e589e41ee69ae5ece4ace5e4e4bce4;
// music[3969] = 256'h2ce552e4b1e390e3bae3a6e45fe4b4e475e6b8e5ace40be6c4e7e9e7ede6a3e6;
// music[3970] = 256'h97e5bee562e7a4e679e52ce573e504e694e5dee48de40be5a4e35ee13ae1b6e1;
// music[3971] = 256'h05e30ae37ee287e3b2e259e18de1e6e2ade305e5f8e705e7e5e546e772e677e6;
// music[3972] = 256'h14e7abe6cde6f3e6f9e68ae66de6c9e611e7efe601e845ea45ea2debb8ecddeb;
// music[3973] = 256'h8feb8beae3e905ea69eafeeb23ebf5eae9eb8eeae6ea03eb9deab8eb6aeb87eb;
// music[3974] = 256'h4fec39eb8cebd2edfbed54eda9ed13ed8dec19ecc6ebcdeb0bea5ce876e87ae8;
// music[3975] = 256'hf1e7aae7bae7bbe75ee880e8aee74de745e78ae86feadeeb43ecc2e83be531e5;
// music[3976] = 256'h3ee5cae65ee90aea5feb17ecf0ebc5eb38eadfea08ebaee99bea19ebcdec94ea;
// music[3977] = 256'h35ed61062d19bc1694163b18e516c015ba15e7177a189318cb18261bc020db20;
// music[3978] = 256'hae1ed21f491f681e891e5b1e891f302184225724cd250a275a28bf29632b3c2c;
// music[3979] = 256'hea2ca52d522d382d392db72cdb2ceb2cb42c2d2dd02c5d2c492c0f2b7c2a3c29;
// music[3980] = 256'h5728f728a7277729f2230412750b2c0daf0b440c760bfa0ac80a880980099007;
// music[3981] = 256'h3e0644069d0534059d049b04e0034e030c03cc02f6022402bd0122019c01c602;
// music[3982] = 256'h320217020200d7fe9ffe1afe2100b6f7a8ebd9eb94ece0ebceecebeb0cec50ec;
// music[3983] = 256'h73ec1ced04ed06ed8bed42ee5beeededdcedaaedccedb1ee14ef33ef43ef1fee;
// music[3984] = 256'hb4ed4eeed1eea6efb2efa1f055f34df499f389f3eaf3ccf3a4f36ff342f366f3;
// music[3985] = 256'hb3f3eaf3d7f35ef4cff422f5c1f5e8f556f874fa7cfb9efef8fef6fddbfeeafe;
// music[3986] = 256'h1aff0bfffafef4fec3fe4eff40ffa1ff8b00b4002b01db014c024a0206029b01;
// music[3987] = 256'h85031507ab07dc066d0691053b0556057a043f027701dc010c028c026c02f301;
// music[3988] = 256'hdf00610028011e01a40138023d02540224026c02c601f2ffa6fed7fedffe50fd;
// music[3989] = 256'h20fd9dfdecfda3fe96febafe14ff70005401ab010703c8021704da0375047813;
// music[3990] = 256'h5e200b1feb1ee41f511d871b481be71bb51ccc1d5f1e781ed91e021f0720d720;
// music[3991] = 256'h03215721d41f091f31204620b4209921e9211022c521bd216621472127225522;
// music[3992] = 256'he2214e212e2149212e21ee213b222a21862039219120b51f3a2117215521b321;
// music[3993] = 256'hba204023191bf709bc061409fe07d508110926091b09d708500921091d09f008;
// music[3994] = 256'hde08d609540a120a0c0aec092d093309160941084708fe073408350913092609;
// music[3995] = 256'hb6092c0ad90a390b3f0b700b510c600cbd0b450cc30c2c0d110d5c0ca80de30f;
// music[3996] = 256'h4f11d40c4504d705ad0bfe0c2111f41318149e15a0143b1349120c10160e470c;
// music[3997] = 256'h580add09f20b890cc10b860c3e0c650c070d0e0d010e760e5f0fc110b7111e12;
// music[3998] = 256'h79124f153d1be12120234022b8236d221f243c25dc2459337841bf4106433345;
// music[3999] = 256'hd045a347c6483e4adb4bed4cca4d714ec64e764e614e4a4edf4db14dd84e7d50;
// music[4000] = 256'h484f944d3b4e9f4e264dbf497846d94455431d427f41af4009404b3f1f3e833d;
// music[4001] = 256'hfe3cae3ba13a0e3a94390739c036d233ec323332ce306930742f6a2eb12da22a;
// music[4002] = 256'hb127b2266526522742275e25eb232c23f61f8b1c351dcb1acb1c042dc535e532;
// music[4003] = 256'h41331832da2e3f2ef52d5e2dfa2c832c162b46292a280128b1270e271c26a623;
// music[4004] = 256'hd7237e1f3b11430be90c520a4209e5086b0750065d0462039e02be01a700fbfe;
// music[4005] = 256'h58fe64fd99fc88fc2cfce6fb75fbe4fa22f9ecf7c6f70ff6bdf58cf4c8f323f5;
// music[4006] = 256'h8de9fed994d872d86ed653d786d657d6ffd5e9d4f8d477d496d45bd4c3d3bcd3;
// music[4007] = 256'h2bd33cd30cd382d24fd2c0d1f4d1e0d1a2d19cd2a4d217d154d099d073d06bd0;
// music[4008] = 256'h50d08bcf46cf5ecfd8cf5dd017d0e5cfdccf64d038d1f5d066d0e7cf51cff5ce;
// music[4009] = 256'h75ce2cce20ce7ace39cf16cfc5cee4ce77ce7dceb7ce78cef4cecece42cef7cf;
// music[4010] = 256'hb4d166d1c3d05dd054d0cdd00dd1b8d0f6cfb5cfdbcf85cf23cf9eceebcf46d3;
// music[4011] = 256'h3bd40ed4e4d4e3d4ccd4b4d48fd474d41ad4cdd4cbd41ad57dd7e9d76dd7b0d7;
// music[4012] = 256'h0bd70fd70ad7cad67dd776d723d7bed628d671d65cd66dd702da5adabdd99bd9;
// music[4013] = 256'h46d898d61cd570d3c7d263d3b9d3d4d3cdd34bd394d399d360d3c0d33ad33bd3;
// music[4014] = 256'hd9d1afce1ace20ce4dce3ccf5acff1cf47d099d017d15dd1e4d1b3d198d1a2d0;
// music[4015] = 256'he0ceafce73cf6fd0e4d03ed29cd24fd2d6d3fcd134d8ece92af01eee20ee4aeb;
// music[4016] = 256'h79ea45ebcaeaf3eb4dec52ec35edf3ecbeecf0ecb8ecf5ec6fedc4ed6eee6dee;
// music[4017] = 256'h55ee66ef86ef1cef8eef55ef57ef67efaaeef6ee8aeff8ef89f057f0f5efeeef;
// music[4018] = 256'h93f01ff1a5f125f2fff1e1f2b5f21bf28cf2cbf1def2b5f3bbf59ff600e962dc;
// music[4019] = 256'ha5dd12de91dd7bde1ede95de73de5ddee4dfa0e153e27fe283e228e254e208e2;
// music[4020] = 256'h7de25de2d1e15ee362e28fe79ff4c7f743f68df7f7f692f74af861f827f979f9;
// music[4021] = 256'h4afa90fa00fbe0fb8dfbc0fb98fcd9fce5fc37fd21fd12fd7dfd06fd01fdcefd;
// music[4022] = 256'hfafd9dfe10ffcffeedfed8fe4afe5bfec9fe21ffceff68ffa7ff3202b1022902;
// music[4023] = 256'hda02e402180370039703c503d40325040904dd04e3066107df0681071b088207;
// music[4024] = 256'hb507f20746078707b1076c073407b0060607e70773080609d40a8b0c2b0b4509;
// music[4025] = 256'h6e0919096d08940827087808ed08bd085a0b5b0cde0b980b31013cf605f796f7;
// music[4026] = 256'haaf544f5c6f4e9f4a8f481f45ff41df4fff456f59df5e8f5a3f437f35af3f5f3;
// music[4027] = 256'h9df3a8f34ef4f5f485f5f3f448f459f47cf4c1f432f507f640f629f606f70bf7;
// music[4028] = 256'he6f5bdf4e2f495f673f61df7e6f8b9f7500017118b14ea1042118a119512f212;
// music[4029] = 256'hc212cf13aa136d1388131814e1142a15631603179c169f16a1166d1639167416;
// music[4030] = 256'h331615162117e817db17fb164b161316d11552166916df156a15f4140a152715;
// music[4031] = 256'h621560156b152416f1151a16f3153515b6158e143a164c150706bffb09fe9efd;
// music[4032] = 256'h99fd7bfea6fd40fec2fd18fee6fe73fed9feb6fe61fe4afe5ffe79fe06fe4cfe;
// music[4033] = 256'h4ffe5dfe79feb8fe73ffd0feb2fea7fe02febbfebffe17ffafff45ff8cff0100;
// music[4034] = 256'h3900d9ff9dff0c004900290197017c014301b500e10032013401de00d900b100;
// music[4035] = 256'h28ffebfee3ff2100da0074010601be00afff05fe98ff10022a02aa021803ed02;
// music[4036] = 256'h0203d4026603d6039004b906e3074c07dc069406d405e8050d06b10519064c06;
// music[4037] = 256'hce06e0072d08c7078c07f407d507c70718083e080509ba080b09e80ad80a080a;
// music[4038] = 256'hd009810931093909790a500b9c0abb093a09e108e508b308a708cc0829072f05;
// music[4039] = 256'h9a041704c503a5038b032a034f032303fe005300f5008d003a001000aa00b900;
// music[4040] = 256'h38001a00d4ffebff82ff8affe000d801db0286044e0481ff56fd6e006902ba04;
// music[4041] = 256'h1907330614054607f506aa046e0fed1bfd1ab919751a2b199718eb18d217ce18;
// music[4042] = 256'ha424fb2d842ce72c402dd12ca92d6a2d352ed42df22c5e3021358c340632c932;
// music[4043] = 256'h5031fb2f9c30f72fa9313933d733c335a0365a38213aea3a153cbc3c663d153e;
// music[4044] = 256'hc03ef83eb43e203ffa3da33d4f3ec33cbb3e773ab7284020aa214f1feb1ea81e;
// music[4045] = 256'h251d9f1dc21cb41bca1ad01928192e185017e515db14ea13df11520fa30d7b0d;
// music[4046] = 256'hd50ca80c3f0c680bdc0a4808a507f907a406e0060c06750517060906eb05fc04;
// music[4047] = 256'he7042404d0033b043b0349055200e8f24def05f12af087f035f086efefefccef;
// music[4048] = 256'h68ef36ef1cef90efc0ef40ef70ef73efa8ef2ff140f240f275f1aef045f0d6ef;
// music[4049] = 256'h46f12af3e9f2bbf20af392f243f2e5f148f1e2f043f0fcef2af037f09af0dff0;
// music[4050] = 256'h8ff09df060f18ff115f1e5f0a8f0ccf00ff1b2f0e2f0aef04af032f2c6f311f3;
// music[4051] = 256'hf6f30ff537f3c6f14cf161f09bf0b2f10df2d2f1d9f251f32df1caee4dede9ec;
// music[4052] = 256'h96ec3bec8beccaeabae8b0e8d7e86fe8dfe7dce7a8e791e7d3e71be775e635e6;
// music[4053] = 256'h7ae694e672e6a1e662e603e762e74ee76be7b6e6f2e66ce61fe634e62ae5e5e5;
// music[4054] = 256'hdae4dde3e4e1c7dfc0ec62faf4f965fac3fb72fb3afcc2fbc4fb64fc4ffda7fd;
// music[4055] = 256'ha5fc67fc15fc02fc7efc4dfcd8fb77fb33fb1dfb69fbb8fbc1fb73fbe8fa76fb;
// music[4056] = 256'hccfb8cfb2efc00fc6bfb48fbb9fa87faf4f98df9f2f97df94ef977f917f802f5;
// music[4057] = 256'hb5f376f571f53ef648f74ff60ef9fcf1bee0dcdcc4de5cdd3cdea8dd54dd72dd;
// music[4058] = 256'h6fdcd1dc77dc16dc33dcafdb66db70db59dbd3da95da02da68d98dd9f0d918db;
// music[4059] = 256'h3edbc4daf9da7fdaf4d98cd913dad5da96daaedad8da5fdbb6dbb0db66dc6bdc;
// music[4060] = 256'h8adcc8dce0dc89dd9cddb4ddafdd65ddb5dde4ddffdd18def0de84e1efe2b9dc;
// music[4061] = 256'hccd4c8d7e6dc03deabe25be54de54de7bfe7a6e761e6cbe310e482e311e129e0;
// music[4062] = 256'h1adf4fde21df2adf87de78df31e1c0e172e2d8e3eae4a4e63ee8dce827e9a1eb;
// music[4063] = 256'h06f2aff434f3e3f39df3e8f347f593f608f917f97b01d911eb17b61acb1e6f1e;
// music[4064] = 256'h9d1fed2021219a22e22209230e23cb2210234c234624eb230c22b721e620541e;
// music[4065] = 256'hf31d9c1ff31e7b1d511d251c2a1bcc1af419081afd19b519af198519301a171a;
// music[4066] = 256'h9d19ee195619d818f118f9189a181b18e0178417cb1770163f15af155f123b10;
// music[4067] = 256'ha20f0b1234204529692690258624a32372239e21eb213821ba1f06206e207520;
// music[4068] = 256'hd61f32204f20951fab1f3c1fd91e7a1ef71d4c1ded1cd61c241c631cd51a8b1a;
// music[4069] = 256'he81aec0f5606fc06c9051205e50481038f036402cd0175012c010a011e00d400;
// music[4070] = 256'h94005f016b0147004702e2f787e724e63de74de698e7cae6cfe6cfe607e647e6;
// music[4071] = 256'h0de636e6c4e621e757e781e765e727e785e745e7a6e7b2e8dee895e909ea43ea;
// music[4072] = 256'hf0ea02eb1beb47eb82ebc0eb8cec8dedc9ed57eea0eea8ee46ef76ef41ef2aef;
// music[4073] = 256'hd5f09bf270f296f298f240f392f450f48bf471f4eff3c9f48cf40af43cf41ff4;
// music[4074] = 256'h96f416f589f531f6b3f6eff61bf76ef9c4fc37fe83fea1fe46ffceffa1ff1400;
// music[4075] = 256'h9100fa00a401dc014402a302c3023a03bb0315045e04c40453056b051a059205;
// music[4076] = 256'hd8057d05340666066b066b07ea07d409960be20ae20ae10a960a4c0c1c0ec60d;
// music[4077] = 256'h870d5b0ebc0d180d110dea0bf30b770cfd0bca0cf40cf30942086009fb08b908;
// music[4078] = 256'h6309fd081d09d108cb082809a7070207b9078208bd08fd08590965082009fc09;
// music[4079] = 256'h29099a0958099f095e0a730a130be10a840bd60ada081208a807d1099e08310c;
// music[4080] = 256'hbb1b8d20421d191fdc1ef11e731fd61ece1fd81fbf1f9e1ffc1f6b20ca1f6420;
// music[4081] = 256'h3c20831fd41fa81f09200420241ff41e091fb41eb31e161f491e601d0f1dce1c;
// music[4082] = 256'h571d7d1d9d1dcb1d411df31c7d1c861c081c571b011c241b641b321c1f1b8e1c;
// music[4083] = 256'hc41b4f1b541c9b105504ae04030523049204d80368038102cb0166029c048806;
// music[4084] = 256'h6a06690640062c062d0663050e0576043e04ef0399031604ab0339041b04f502;
// music[4085] = 256'hff026d02a103df02f6034110a117be152d1688158314d814201438140a146e13;
// music[4086] = 256'h1c1380125c1284123a12d211d21198117f11f711941132114611dd10ba106910;
// music[4087] = 256'h6c0f630f7d0f180fa6101b121c12b81356140813c2125a12e311b211ee108510;
// music[4088] = 256'hbf10a410d20f690f130f6c0eac0ee10e1b0f910f130f8f0e5f0ec10d250d520d;
// music[4089] = 256'h050d740cf10d190e580cf30b230a330856088c0711073f077a07ec08ee088e07;
// music[4090] = 256'h1f07a40617068605e1047b0400046803d600ecffa90142f9c6eb1be9bbe975e8;
// music[4091] = 256'he2e861e836e883e8d7e7a8e7b4e7dfe7bee7c6e787e71ce7b5e72ce720e78de7;
// music[4092] = 256'h89e6e0e6e4e65ae6f6e536e4c1e394e492e546e57be5a0e633e42eea74f886fb;
// music[4093] = 256'h7cf987f99df8e8f9dcf9ddf878f945f9acf9fff937facbfab6fae3faadfaa1fa;
// music[4094] = 256'ha4faacf92cf942f93df93df949fa95fb4cfb30fa9af8b5f776f768f73df851f8;
// music[4095] = 256'h6ff839f8aaf73af9d3f990f936f948f82ff8b7f694f6a1f67ef507f7baf564f6;
// music[4096] = 256'h6cf6a8e8f7de6de022e068e08ee07ddfaddf93dfb2dfd0df3ee012e0a2dfe1df;
// music[4097] = 256'h3ddf74dfacdf4bdfefdfc5dfb3df47e092e0d9e0c0e0a7e0b6e042e178e14ee1;
// music[4098] = 256'h91e116e125e1a4e194e116e257e294e272e2d2e1bbe165e171e1b3e1a4e1b0e1;
// music[4099] = 256'h1ae116e1abe1d8e127e23ee203e21ae281e2cae266e3d1e38be2dde1c7e2d7e2;
// music[4100] = 256'h67e3cde568e79be787e738e717e810eadaea07ea7de8e7e74be856e886e801e9;
// music[4101] = 256'h04e982e841e867e89be81fe912e9ace8e7e810e967e9a8e96fe92bead9eb1bec;
// music[4102] = 256'he8eaa7eabcea9fea10ebf1eaceead8eaedea57eb0eeb29eb44ec37edf1ecdaeb;
// music[4103] = 256'hfcebc1eb4cebbaeb3aea7de8b9e8eee805e9c1e943e9fee681e6e3e64de6c2e6;
// music[4104] = 256'hb5e6b0e646e7bbe624e7a8e7a1e7fbe78de7cce707e8b8e7c9e713e7e6e694e6;
// music[4105] = 256'hebe4c4e3d4e322e557e501e666e94aeb97ea83e53ee29bee97fe850363055706;
// music[4106] = 256'h2205530588053005eb04190450031103ac023002f501c700c000af0096ff7c07;
// music[4107] = 256'hd41229146113de14ef14d9153316bd14da14c4190b1fd71d9e1bbc1b071a3f19;
// music[4108] = 256'h381a871a311c751e20207122c72313255b272d283c2a6f2c3a2c592f692dc11f;
// music[4109] = 256'hb818b51ad519d319511a3a19e5190a19cb17a217a015d514be14a613cd139e13;
// music[4110] = 256'hf5125112df10c30fc80e180e920daf0c390c280b6e0a8f0aa8086a06ad051505;
// music[4111] = 256'hb20448043e044c04f5026901a9004300a0ff92ffbf00c1006b009b00ceffceff;
// music[4112] = 256'ha3ff89ff9300d8ff46019a00d0f596ee52f072f041f062f1f7f00af1bbf25ef4;
// music[4113] = 256'h82f47ef409f51df572f5fff4bef4a0f646f7c6f6b8f6b2f57af519f6ccf59cf5;
// music[4114] = 256'ha5f598f579f55af562f553f57cf5a1f5b4f615f9aef9eff8cef850f830f877f8;
// music[4115] = 256'h39f83af8b3f87df91dfa63fa5ffafff970fadefa41fbd8fd2100220073ff36fe;
// music[4116] = 256'h5dfd7bfc93fa53fa71fb7dfba7fb0bfcbffb28fc2bfc71fa08faf5fa73fb28fd;
// music[4117] = 256'h6cfeeafd39fea3fea0fee5fe8efe76feaefef5feb8ffcefe9bfc55fc7ffd11fe;
// music[4118] = 256'hcbfe03002e009100fb002e00fd00fdff35ff5b0a7b165c166d15dc167f15ba14;
// music[4119] = 256'hfe14d315f9162a17a017a417ac173f1813188f18cd18ea18931adb1a881a5c1b;
// music[4120] = 256'h3a1bf81ac11a231a241a451a6e1a7c1ad61a901b901b271cb31c741c071d321d;
// music[4121] = 256'hbb1d491ed71cd21c851d541d181e011ede1e0c20f01f6822201dfc0d9508e60a;
// music[4122] = 256'he509080a5e0ad309b30ae6092208690720072307e0061a075f072d07b807d607;
// music[4123] = 256'hbb071e08d80797077707310759079b071d087b085c083708450817095d097808;
// music[4124] = 256'h55085b080b080808df07fe071608c107cd073f08f0086609a9090d0a290a4a0a;
// music[4125] = 256'h270ac209d309cd09db09e409c009df09ef095e0a010b650eee11700a8c022208;
// music[4126] = 256'hab0c870d771213146d14a415d01369145a149010bf0e870cd809b60894065b05;
// music[4127] = 256'h86053a05d8043805780743096609320a3d0b450c920d8c0ec00f0b1387183a1a;
// music[4128] = 256'h45187419fe190e191c1b9f1b961cfc1f422070266a35ad3c4f3cbe3e8840753f;
// music[4129] = 256'h7f3f7d402241a6414a42f6425043ab43a04317438c426f40d13d0b3ef93fbe40;
// music[4130] = 256'h6a3f713d5d3cfc3ad839bc396d382536e13407356235fa3463340e3312322a32;
// music[4131] = 256'h1131c13059304a2e3d2ee82bad2bc3379440a03de63b593bc738f43612379339;
// music[4132] = 256'hd338be3578356333b330c82f012d212bd22a292a022a3b29ed28c028ab277727;
// music[4133] = 256'h7a26a2254a2571226520a41f5d1eed1d681c151bab1a881960196f175416fb17;
// music[4134] = 256'hb710c2047601c50187008fff4dffbafe96fe49fffff626e852e425e658e490e4;
// music[4135] = 256'h7ee4fce2dce2c9e1e6e05fe026df7adec4dd53ddcfdc44dcb4dc4fdc7ddbe9da;
// music[4136] = 256'he0d9d0d90cdae1d9d6d99ed9d8d9c3d934d9e8d866d866d853d8ded7a9d7d9d6;
// music[4137] = 256'hb5d633d75bd72fd80fd854d74cd764d6e1d530d646d69fd666d620d656d670d6;
// music[4138] = 256'hc8d60ed764d746d7efd6b8d7f9d719d8a1d817d933dc9fdeafdd0ede62de86dd;
// music[4139] = 256'hd2ddc1dd77dd25dd97dcc4dc68dcf3dce8de38dfa9de3ddededd04de09de2bdf;
// music[4140] = 256'he6e0b7e08ce05ae148e1d1e0d7e010e192e14ee28be29fe212e33be39ae339e4;
// music[4141] = 256'hf6e3eee335e4dbe34de4d7e4ede4b8e664e8d6e714e7ade666e6d6e548e49ae3;
// music[4142] = 256'h83e3a5e2cfe266e35ce388e38ee3cce354e34de231e3d9e290e0b5e081e1b0e1;
// music[4143] = 256'h10e314e486e391e251e3b9e443e447e430e56ee5dbe579e534e575e5e2e485e5;
// music[4144] = 256'h0ce574e3e8e334e286e5e2f3fafb5dfa15fbf6fb9bfa26f944f8dbf90ffbddfa;
// music[4145] = 256'h8efb79fb78fb50fc78fcd8fcdcfcadfc33fde6fc70fc97fcd0fc00fd7efc19fc;
// music[4146] = 256'hf7fb86fb7afb44fb56fbccfbaffb4afccffca2fc4cfd84fd16fde1fcdffc2efd;
// music[4147] = 256'h19fd89fdfbfd13fe18ff48fef3fe9100bbf6a1ea82eae3eb11eb05ec84ebebeb;
// music[4148] = 256'hd7ecc9eb3cecccec0dec17ec2eec26ec4fec41ec53ec54ed8aee0fee51ee01f0;
// music[4149] = 256'hf5effbef27f03eef02f0c9f008f144f215f260f222f4a4f48ef4fbf3def3f7f3;
// music[4150] = 256'h14f33ff4f7f335f3fafbaf0531068705fe058205d20596056a05140631066e06;
// music[4151] = 256'h3f068d051306ea06120754077907a1074209ce0a8d0a1b0b570c150cf90b1f0c;
// music[4152] = 256'had0bf10b790c110ca00bde0b980b780bcc0cf60cab0c4f0ec20e050ebe0d030d;
// music[4153] = 256'h830d390e9b0dba0de20de00d550eef0dcc0d590e780e820e4c0e500eef0e060f;
// music[4154] = 256'h8b0ee90dd70ce20ba70cc10ea70fff0e940ec70e6d0e560dac0bf809d909ed09;
// music[4155] = 256'h8009150ac0084b07cf0843082708d409d008890a2d093bfd31f67ef66cf45af4;
// music[4156] = 256'haef53cf5c9f5b3f5acf5ecf60df74bf7cff749f740f75df74af7b4f77af778f7;
// music[4157] = 256'h8ef6ecf3c5f945089f0e1a0d3d0ecb0e2d0da00c940cc90c7e0ccb0b9b0b2f0b;
// music[4158] = 256'h820b010d120e110ed70d380e530e310e5f0ed80e231006108d0e560ebc0d0f0d;
// music[4159] = 256'h020d8a0c930d730ec40d840dfe0c6a0d6d0e220e780eae0eda0e600fdb0e870f;
// music[4160] = 256'hd20fc60f23114f10801263133d0686fb11fd8ffc8dfb9cfca3fb4bfcb5fcfefb;
// music[4161] = 256'hb4fc19fc8cfba5fb92fa5cfa86faccfa7afb45fb96fbdefb54fb83fba4fbe0fb;
// music[4162] = 256'h60fc12fcf6fb16fc12fc3dfc1ffc1afc33fc16fcd7fba8fbf6fbe4fbc7fb26fc;
// music[4163] = 256'h53fb7afabcfae6fa57fb40fbf3facbfb01fc0afcadfc60fc38fcdcfce2fcaefb;
// music[4164] = 256'hb4fa6efba0fb6efbe3fc5cfd7efd97ff1701d00125024e017f014d02f001d901;
// music[4165] = 256'hf901350165000600f5ff31002d0097007402e10378030d03e902010135feb6fe;
// music[4166] = 256'h16035f06e905a5041e059606e8068204fb02b407450d7e0ce509ce07c8039600;
// music[4167] = 256'h13fea5fa2bfb7901230681015ef539ebd6ebb9f3fdf272e550db16e4b9f99a04;
// music[4168] = 256'hbe00e7011c0d3b156e0c12f84cf1fdf843f92eea5ad109c27ececfec3d05910d;
// music[4169] = 256'hd20c1b0aab0718086c076705350768080907fc0937136a17f90ddf050a0c9b19;
// music[4170] = 256'h2f22021ae7086104e110c21e0e1866ff6de872dd2df0511c2b40b8520451413a;
// music[4171] = 256'h8d25311dbc226e37ec454c3d2724480c5205b50b5313011a5b1f3c1f021e8624;
// music[4172] = 256'h122cf128f01e2b1c1b25fc2afb26d4232a2693318641ff422e38312f0a286324;
// music[4173] = 256'h892468263b30373fdc4a3456b65bbb511247e0464148d54c1b54e156e0603e70;
// music[4174] = 256'h446d0e5ce452a059f06a2a77af76356cd055d83eff323a2853191c0440e979dd;
// music[4175] = 256'hf8e1c1de49d931e7a9fc130113f5c4e140d0bfcf29d86cd838da67dfd5dd5edc;
// music[4176] = 256'hb2e1faed4bfb4f03060d7c1588167319ff1f33283431c834583484344f37d237;
// music[4177] = 256'h4a2a601958195320971e25199515cd12b314e81cdc213c1de3146212bb17a41b;
// music[4178] = 256'h5a163f0d990cee1227183321d028e6205f0922ef55e60dec41f33afe170460ff;
// music[4179] = 256'h83fb0203b9181d2e9636bb35e32eb92190126d0482f5b3eaf2df9bc93ebd77d6;
// music[4180] = 256'he602d51fb125c021f1267f31ec2b721e091c6924802b7925a11d53206428302b;
// music[4181] = 256'hd820a514281180132b187a16060f720d0819a12a01324c31e230e72eec306937;
// music[4182] = 256'h1d36202c0a26ac2e98407d4902494b4d13535e502348773fcd3eb1487b4b3e46;
// music[4183] = 256'h3e45f2477b5552604a5d8765a3717d72e96bb2542d3e9a36ad2e71230516b610;
// music[4184] = 256'hcf15a3148d18d924fb289e2dfc2c2d2002235738d2483c4a584244406a441b46;
// music[4185] = 256'hd7450744063c5d2fcc2b46308a2c371f0417741dc3238c1e4515d30c3b0d3615;
// music[4186] = 256'hf11d4d2a41265e08dcf662fb3afb39f6dff3fdfad407fc06b306f70522f068e4;
// music[4187] = 256'h7bf7fd17b82d0f2a02217324bb2dd031b82e962b5a2cc035c84132490948dc38;
// music[4188] = 256'h9e27b81bdb15ea1d18311a430a4bf14f2055d85a935731378116e9149c1f6f26;
// music[4189] = 256'h882c5838dd3ee939fa333e324b356f3339321939f13768305130243cc4443e3e;
// music[4190] = 256'h403b2b40584054382931f734d43b95416144b33ee0395b37c932a136a93c4b34;
// music[4191] = 256'hc02cba2ca42c6d32cf2aa5121a0dd619112404222a0eaff366eed105271d3c1e;
// music[4192] = 256'ha90af7f294f2090ba31b75114cfa2fe49de4b5057e1b95141911ea126e135a17;
// music[4193] = 256'h3b16d80fa1121e1cd31e6f1b60132f08510aa518021a3111fa0a51f78fe3bce7;
// music[4194] = 256'hf4e94ce70cf616051a0724fc44e58cdbbde4cee9b7e1cad519e215001908af02;
// music[4195] = 256'hbb029506cf073a01aa1011330d3f103c3a325a2051196d1b6d21b22a882a4f24;
// music[4196] = 256'hb1208e1bb118241a991fb7293f25830e91038a0f5919f810310c79165e203423;
// music[4197] = 256'he71bd113521a9d26b729771ff413c21818299f31102aa421e62405203e072df6;
// music[4198] = 256'hd501901bd72c7e2af616b4074b09ed0e7514ab171416101b2f1cc715ea15860e;
// music[4199] = 256'hd2fc62f043ed96ec85ea17ffdd1ed422501acb13550bca097f10451bc81ce812;
// music[4200] = 256'hc20aaa09f612d5113301a5fe72f717de8cd2a8d52fd907d729d884ea42f993fd;
// music[4201] = 256'h6601aa0025fefff74ff280efcaecd3f287ef36dd59d630daa6dbe2d6c5ce35ca;
// music[4202] = 256'h64ce48e104f495f26ceafdeddbf483f53ff053e581dd43de11e0bae30eed41ea;
// music[4203] = 256'h7fd1d9c251d1f8ea5cfc7af7bbe292d4f7db97f04dfae7fa96fb1dfadff712f7;
// music[4204] = 256'hfef929ee1dd6bad06ed0cccc92cf9ece06cf9cd0a6ce84cae5c679d82aefcef4;
// music[4205] = 256'hedf794f33aeed1edede7f6e617e4e1e328e68fd024be19be81bad7b8b9bb32c1;
// music[4206] = 256'h56c062b47eac4bb0f4ca88ed46f130e1b7d954d785ce9fbed2b302bae4c54dc9;
// music[4207] = 256'h02d4a0eca5f62dee56ef79f6dfeba9d6d4d22ee6e2f40cf49ef8830597073dfd;
// music[4208] = 256'h4af91af651e517da47e53efc660436fa48f7eeff2f0be4100810c706f3efa5e6;
// music[4209] = 256'h75f55a08391054fd73e40ee12bec13f240f221044a19e91bc819d917071159f7;
// music[4210] = 256'h37daaed76fdaa0d58ae025fcf10cc105a4fb31fe9f001ff41ae547e590e979e4;
// music[4211] = 256'h0ee69af88e04beff24fdf20007f8b3df57d52ddbd0deb6e184e1e0dd0edb8ee5;
// music[4212] = 256'h1cfe1202bfec53d570ce0ce0ecf2b8f4ade42eccaac1a7d2abeda8ee0bd848c4;
// music[4213] = 256'haec170d4a8e423dd59c6b3b9b8c218d39adde7d31fbd50b2b0b910cfdad8d4cc;
// music[4214] = 256'ha3ba22afe2bc53d5d6dd61daa7d705dc37d153bb49b95abbd6b8c6ba31baf9ba;
// music[4215] = 256'hf7bcb8bd7dbebabce3be41c13ebfc3bfbebf0abf00bfe4bd0cbd2abb30bdccc1;
// music[4216] = 256'h7dc2b1c282c02abd98bae2b426b7bdc36bc90eca0ccdd4cdb3cbe1c5ccc956dd;
// music[4217] = 256'h20e409d802c677bc76cea5e5e9e608e15ce28be3fadd0edc04df86e0dbe2eee2;
// music[4218] = 256'hd2e115e3ebe229e133dd3ed79dd403d954e855ffbf08d6030afff8f6b2f283f3;
// music[4219] = 256'h39f353f996ff09058d045bfdcc02fffbf2ddb6d1a7d723dbdddc16df2cde01db;
// music[4220] = 256'hdde7f7fdbf02e904500e2d13dd15bc12af0a4e0564046608f9077305c406f209;
// music[4221] = 256'h1f0cbe0b000d0d0a8e0be811e3066efbc8f41bedf6edbcf2dffb50f737e9d4ec;
// music[4222] = 256'hefe6a9ce49c397d298e93eee50eb22f404fd7ceac0ca62c883e2bdf9bbfa0bf7;
// music[4223] = 256'hdbfa77fac1fb51fcc7fda9055c09d308e10266fed4014803f004630a030fd10d;
// music[4224] = 256'h7f0deb10f612831531154a150316ea14dc17bd0d9bf8e9f25ff9d5f9bbf5bbfe;
// music[4225] = 256'h78140d1dc40b76f585ee23f137f23bf38f07b5208b225421d125a12874297e23;
// music[4226] = 256'hfb220e27e425d121d0209025e025a2238627c229aa245f23a22ad42b262bf728;
// music[4227] = 256'h3e24fe29ca24c10b9ffb46042c1e932d19221709c200ef09190ba9081613f42a;
// music[4228] = 256'h5135b620e9077f0180139228672b962b632a4225f42301237c24be2863264021;
// music[4229] = 256'h5b2284237324c5259123c121a71b1d1aa41d911bcf1db51a75127e1260122f11;
// music[4230] = 256'h690f4812f311b90cd118f72d0a35d822b20e7c106d11b30ddf052dfc39f9faf6;
// music[4231] = 256'he20900224d210a1faf1b3117be197a18f917131dcf2214241220d0177b0e0c0f;
// music[4232] = 256'h3d1479104708ff084f06e5ee39e3beedd6efa9ec9be93ceaeceffade74c12fbd;
// music[4233] = 256'h13ca68ccd6c815d385e016e239e218e68be236d1fbbe7bbe86d251e41ee0fdd8;
// music[4234] = 256'h97db2ce061e3f3dd82d893d9fed9dadb69dad7dafcdc03d774d5eacd90b8f9af;
// music[4235] = 256'h40b1eeae08af69bac1d1abda49c509aaaaa557be87d86bd9ddc065a21da1c8bd;
// music[4236] = 256'habd959dd9ac117aaeba87da9a0a70eac5ec349d56fce64ccf7ccb0cae3cb7aca;
// music[4237] = 256'he0cb83c94dc5adc701cd27d71ed398b772a42aafd7c5a2d287cb67b2dda633a8;
// music[4238] = 256'hb6a05aa59bb4d5bbe6bea6bfb4bc13b39dae40b5a8bb63beb2b7a5b0d6c14dde;
// music[4239] = 256'h83e285ceeab9cdb9eed12eddefd490d8e1e077e307e2c1e091e614e974ea9ae1;
// music[4240] = 256'h7fc72fbf68c689c495c033bea1c0aec6f2d3c9ee75fb15f6b6fad806b50dd90a;
// music[4241] = 256'ha8086f0f6016101b861698115812ba0094ed9ceb9bebe4ec6feefeef22efb1f1;
// music[4242] = 256'h7f09771f8d218c216d21ef1b931a7022e71fb40877fd1213fd2c1c32712f7333;
// music[4243] = 256'h4437f42a7f1069080917a81c711ce21fb81af416b319a11ba920472212250d27;
// music[4244] = 256'h9d1258fb76ffc218602986231821df28f6264b15ce003bfdf70bbd1f5e231620;
// music[4245] = 256'hc02dab2c541352055a047703480029073b1bad1f0a08aeeefae84fee87eb8fe4;
// music[4246] = 256'h1ef2f60917116212fc10830aeb09e1122a1ca60b9df161f0d3f429f47bfa3310;
// music[4247] = 256'hf12ae42cd417ba07f107560cb00bfe15d72fb33fec338b194908341465373a4e;
// music[4248] = 256'h0d45e1296a17a4153e19311f542c45418c47f337ab296228333b2a50a34fdf48;
// music[4249] = 256'h1d4a144cc73b4628b32eab44c4591257d53a5d277a27f12b4927872a93416653;
// music[4250] = 256'h514dc1361b2e6f33b9309f2db02f72346434e42d4929e421f127ae43e3535447;
// music[4251] = 256'haf33a5290026ba2f2a3e9f408b40013f6f49c36042635151df3f723ba73ee83d;
// music[4252] = 256'h403ece37a72e23362e4f3366c65a893a4a29232a8a2f262ace2d92451454d655;
// music[4253] = 256'h0a552d55ed51874bec4a1a3fcc27bb21c32bc82b6e244631323a03284a1e1e27;
// music[4254] = 256'h5b2b471b1502a5fb1401b5fd3cfa4107b01639175917591ebf1ce607d5f3dbf0;
// music[4255] = 256'h6aedb7e87af179075f17140c88f46fe8d0f2af08d0111e1116113a133e0cc1f5;
// music[4256] = 256'h28e992f01ffff2047dfbafee05e926f3ca03f00104ed9ed9f5ddcdf7ad0bd605;
// music[4257] = 256'h34ee7cdbeddc89f05802aa0121ec9cd497d55ae8a6fbadfc9ce66bd727d6add7;
// music[4258] = 256'ha0d763d551d402cd38cf07e8a4fbf3f5e2e184da81dae5d027cdc1d1f2d69dd9;
// music[4259] = 256'h3bd3d2cbfbcc72d58add90e060dda7d499ce8ccd95cde7d081dbc1e74cea9ae7;
// music[4260] = 256'h13e416ddbdd956daaade16e507e2e7e41bfa76080907ed041d066eff8eee12e6;
// music[4261] = 256'h2de901e8ace181e668fb940af80bcc11e21d35208519531a7c214a28322ee12a;
// music[4262] = 256'h60213e1e6c24732b692bc5277320c11b3c1f8723bf2a08321d320e2dd527f029;
// music[4263] = 256'h9c2560106b039f0ec52482303922ca06fafb7709671f902a832366104d05a412;
// music[4264] = 256'h621bce116011681334137217bf163d170a13b007b403f206ff092d041a014207;
// music[4265] = 256'hb20b380e0806a0faa4f611f184eef2f0edf765f41adc41cc8ec8e9c584cb3ed1;
// music[4266] = 256'hc3d1c2cf6fcb84c9e5ccc6d299d680d4b9d037cd57ca03dbf7f543f829ed32e8;
// music[4267] = 256'h53ec0cf424f31bf3e7f32ced03e650e16ae5afec08eb7ee56be302e782ef08f5;
// music[4268] = 256'he1f0dcec1de7f5d6c9ceafd808ebe3f1baeb67ec8aee85f045f39af13bf094e9;
// music[4269] = 256'hd2e464e4c2e440e97bddb4c5afbca5c94ddbf0dc27df8fe775e773e5e1e3c3e1;
// music[4270] = 256'h07e18ee08ddd1fd890d417d6f4d9ebdb02de6fdfe9e0a1d738bb87ad4eb3e1b6;
// music[4271] = 256'hb8b5a3b8d4cdafd956d62fdb57d8a3ddd8f036f92af7d1f274f3c6e6d9ce87c9;
// music[4272] = 256'h4ad18ed86adaa6e74afb4cfae3f7a1fb34fc96fe49fc4cfa66ffaf027100ddff;
// music[4273] = 256'h8105c909480a9a10a31041f845e37ae8eaf9d10566ffddf3ceef4efcf4121c06;
// music[4274] = 256'hc4eb1df01afa1efb50f755f180e7bbd983daf6e910f804f45adfe3d023d254e5;
// music[4275] = 256'h39f9d2fa77fa10fe12ff51fe8ef8d1f263f216f752fffbfe0cfc60f652de9dd0;
// music[4276] = 256'h3bd6bed41bd4cad551d99be076e33be24bd748d98bf15af910f359f57dffdffc;
// music[4277] = 256'h9de7e7d95acfaec77ed117db75dc32d786d088cb14ca0bdf7bf634fa0ffcfcfc;
// music[4278] = 256'h65fb4efbd9fa8ff793f13af47ff387e04dcebdd4a9eec0f9c1f520f4d3ed2ce7;
// music[4279] = 256'h22e848f3cef3e5d866c3e1c67dde22f06de53ed482cdc6db4af196eea9e698eb;
// music[4280] = 256'h76ef2ae9bce5f2e63edca7cc3fcbeade03f01bed43e8c3e432e534e8e5edadec;
// music[4281] = 256'h6dd1c3b983b497c2d4def0ea97fd670e8307860a1a137a083eed2ce136e705e4;
// music[4282] = 256'h2ae21ce645edb3ee52eab7ecf7e81cf31009a70cf0087304e7ffd7edb1d981e0;
// music[4283] = 256'hc0e802e643e420f29105e00505049a044101d9f50cdbdacf0adf8bee1ee7bdcd;
// music[4284] = 256'hd7c19dcff7ebc5fabdeb60d155c207cfece665eee0ed24f19ff17deccdea7deb;
// music[4285] = 256'h17dd94c8eeca40dfc1ed62ecd2daefc8a9c64fd504e877eb42dde1c8e4c34bd5;
// music[4286] = 256'h57e763ea15d7dac330c56ec64fc72dc8f9c20dc4b8c4fac840d09acad6c49abe;
// music[4287] = 256'h9cb97ec090c3d5cbe3dd02e48ae379e5efe665da92c11ab957b961b99bc4d9cc;
// music[4288] = 256'h01cd0cca98c2e7bc85ba38bd53c5f0cb94cef2cdacc8c5c3a5c131c893e081ef;
// music[4289] = 256'h27e737e2aae424ed6ef345f003f033f0cdf2f1f30aed39ecdce65fd5bccb06d6;
// music[4290] = 256'h7aecadf89bed86d744d047e224f819f90ff481f95df9d6ff1b103112180ff20c;
// music[4291] = 256'h830efe138512df0e790faf1afc1d4607d1ece0e362f5940dbe1a10228f1eb313;
// music[4292] = 256'hb507a0069b13511c9b209913cef7a2f06bf6f9f51bf6f9f548f40af3a8f62800;
// music[4293] = 256'h7dfd0ef96c06590a2c0600088a09ad0f8510a90e5e0e590c2b10a20dd9117316;
// music[4294] = 256'h450200f155ec74e883e2aae760033d14d11361136f111b0e6d10751b2f1579f5;
// music[4295] = 256'h72e114ee22074410c111cd160018eb12e110d11388080cf283e70cf4f1062b08;
// music[4296] = 256'h90094a0e730e440ffb08df05ae066a0a7d0ddafa84e821ede303d7152f0bb9f3;
// music[4297] = 256'ha0e3b1eb03040711cf10330c1f0c3b032bee80e327e1d1df7be1d1f1e6072d0b;
// music[4298] = 256'he7040306290adafecceceeea23ec3fe738e639f79e09c7084808c1090807cf04;
// music[4299] = 256'h5b060f0802f2ffdcfae190e841eb40e8f4dec4d9fcdb7fe0f3dc64dd05f12e10;
// music[4300] = 256'ha81a6f057cfaed06c31395168c083df367eae1f8f413571e9e0eeef5cdeaeff6;
// music[4301] = 256'hbb0abf10e80422f2faed0602d7165f1a03169e11c6078bf626ea06eea0003111;
// music[4302] = 256'h031242106e107d037ef5bbf596eea6db7cd718da0dd266cbb0c9d9cc59d754dd;
// music[4303] = 256'hb7de7fe13fdd7fd8efe1ecef30f5caefe9e223dae1dd5be917ef9ce9b5e094d7;
// music[4304] = 256'h11da61f4300c010972f78de9bae6cee237d611dce4fa1b0e5f0690fd64031e05;
// music[4305] = 256'ha4f417e388ea9503340dd506e7049b08a5071a025002b501c1fc76ff44048d05;
// music[4306] = 256'h1d08d90a6b094a0291fbc7fb680034012903850382f041dedadf1ae0a1d7dfd9;
// music[4307] = 256'h78f3380a690382eb8ed7e2d8b1f0c608bb0d8e003eef96e425e542e835f37a08;
// music[4308] = 256'h3c0dad0a05110813931392136a14e3131d103e18831d4918b31834152c18b22a;
// music[4309] = 256'hcd3146301a2ca8146201be0d67283a3b9933b60c04f38dffcf097506f907f905;
// music[4310] = 256'h5807730f550f130af70a1a1ce82a9d1f6c09e3f903fe710c7d0b9807980ad80c;
// music[4311] = 256'ha3149a114ffdf5f7fdfc53fc8ffea4fec6004a0373035105d2f4b3e621eee9f2;
// music[4312] = 256'he6f5ccf757fbaaf9eef2b2074c1d501e462124246629ba2f0e34b62b790f6703;
// music[4313] = 256'hc50af3137c1c5b1b2916060e95163736453f7e380a39b236df374c39f239c63e;
// music[4314] = 256'ha442ac46bd434940a140d830581d0b206233713f023be53a254672438d284910;
// music[4315] = 256'hb3152c2fa23d7c371c3265372b358720ba0f121aba2f4a39d4369835db365a2a;
// music[4316] = 256'h7d14a60a7718952e4c33583080306532c435f4332d31d82b252b9c2ec3189200;
// music[4317] = 256'h4e05f50ea30c560a17163e246f1f2c12230dcf0b760f87173c1c6b2f00485b44;
// music[4318] = 256'h722e821fb91d28198d102e1c7a377c467836831bd10edc0e881550198a28ac3c;
// music[4319] = 256'hf736d12e9a309133e936dd38403b94295710050dd0180e32aa34960e23f4d6ef;
// music[4320] = 256'hc2eae4e9a9f6b311b625e918e8f9bae987edb7f2e1f085f9e0106d1c410efcf8;
// music[4321] = 256'he2f2fbf69df6e8f5fa04a01df31f810aeef22ce94cf961112a2089285c2d702b;
// music[4322] = 256'h2e1474fb43fa53fc7efa36fb45fd15ffad01850e361b701648054bf775f8fbfb;
// music[4323] = 256'hd8f8f2ff6f13e81ed61382ffe6f8f6fba1f812f181f7470f381e6f13f100b8fb;
// music[4324] = 256'h47fe20fae2f03fef21f4faf697029813591470066bf496f80219592c6e2ca728;
// music[4325] = 256'h66257e21e10e3e03b60c281111091602d811e12a752c1e1ae60678ffa6fb84fb;
// music[4326] = 256'hef0a58231a3e9841bf27a617921d8523c922ba2fdd419d3e2636243c6745f336;
// music[4327] = 256'h5b1e3e1a5f1b501a371b7d1db01f2c1cb0274e3b7a3a33286915cc1c2f361144;
// music[4328] = 256'h973ac41db70eb1081ef76df270006b18fe28151936feb2f6edfac6f921f8f006;
// music[4329] = 256'h891ed4276919d10087f83809aa218226f0106bf702ef29fe3c13bc1dcc266c2c;
// music[4330] = 256'h2227980d24e608d7e7d9dbd79bd804dba7e1a3e983eb7ce6aee0e0f0fd06a206;
// music[4331] = 256'heff91eee40e968e035d68ee51c0603172205e3e373d689d818d8eedaace5ffe9;
// music[4332] = 256'h00e122d898d522d5a4d514d362d019df52f6d3f85ee721d401d17be254f17cf3;
// music[4333] = 256'h5bf589f88bf712f5aff263e6ffcfafc736d0bbce1ac507cbf8e265f3c6e3d2ca;
// music[4334] = 256'h85c2d5c15ebe99b87fc07cd374e61afecf0442fc3df4a1e360dd6fe450ee40f7;
// music[4335] = 256'h37e558c8f6bbf1b9edc07bc718c9c5c411c26fd416e661e600e5eae14ad830c6;
// music[4336] = 256'h9ab9c7c253d63de085d2c5bff5b3a7a02e984f9e56ac92c87ed118bf9caac6a0;
// music[4337] = 256'h67ae38c395cd07d2e5d321d3b0c95dc305c4acb868a7b1a6d7bc36d1c1cf09c8;
// music[4338] = 256'h32c94dc946b6f1a01fa9a8c7bde168df0fc618b3e7ad54b062b45ab588b365b2;
// music[4339] = 256'h05bc1cd0f9db18cf97b601aee2b344b878b808ba87bcfbbfb9d19ee7d3e994e4;
// music[4340] = 256'h1ce81aea13db55c5a1bfd7c123bf04c2a9d4c3ed0df251dfb2d2aed47dd3d9c8;
// music[4341] = 256'h8ec6cfce73cfeed1a0e10dec23ec31f185f812ef3ad770c989cacfcac8c775d1;
// music[4342] = 256'ha0e9f5f7b4f62ef770f75ce46bc4e3c78ff46f143f19c0072ce9a6e2b1f4690b;
// music[4343] = 256'h3a16660698f40af036ed78e919eb44feb712551462135716ad108bfd2fed50f5;
// music[4344] = 256'ha709bf120b0d4ffbfbefc6fcee092200ddec41dbdbd47fe58efde705def685e0;
// music[4345] = 256'hedddaee3b7e096e01be362e474e236de2ce0acdfe6ddf1dedee090f193014bfd;
// music[4346] = 256'h65ee63e056e686fbc70705027af122ee88f717f858f350f364f501f689f525f5;
// music[4347] = 256'hd0f617f335eb0dec26f21af842f82af483eee4e502fa151bf71ce7175314650f;
// music[4348] = 256'h3212c213141cb520c31b8a184f07bbf8d5faf9f7a2f4f9f28ff023f4d7f719f9;
// music[4349] = 256'h23f114edaa044f17c214e415e2166715b813c412b7141e0e8c092f0cc70d8112;
// music[4350] = 256'h0410b10e2a11c8fe20ede6f89e123b25b82a5b29fa2687279a2d4a346b305418;
// music[4351] = 256'h6cf996f5cd0d611ece1df11d4a228423f122f824291e300840f22df113083916;
// music[4352] = 256'hd11079118810cd01b3f5c3f234efffebb4f030f5b3f82bfaf2e78ccf9dcbf7d3;
// music[4353] = 256'ha6d44bd185db49ecf0f162f3bff8e4f4f4df25cb82c814d1fdd429dbe4eb1bf6;
// music[4354] = 256'ha7f155ed1df31ef419e200d1a6d1e5d646d536d8b8e8c9f3fff4adf85bf945f7;
// music[4355] = 256'hbef733f829f52befacecdae669da8cd66ee366f768fc5cebb9d625d414e700f8;
// music[4356] = 256'h82f63deaaadeb1e08af29cff87f767e717e14ce7abf7270204f844e426dad7e5;
// music[4357] = 256'h6efe520849fa76e2c5d13fdca5fac4093a0b2c0ae6fd8df368f3bafb1805c3fc;
// music[4358] = 256'hb3f133f0a3efb8f671fc04f9dff47df1b8f3b4f658f25dee2eecd8e94cec0ef3;
// music[4359] = 256'hf2fa8000b2feb3f86cf32ff14bf1bef01ef5d7fb51ff2000f3f138dcabd32dd0;
// music[4360] = 256'h23cfb2df5bfab504c2fe39fa9df6fdeba0da56d42fe5d9f89afff7fc84f771f4;
// music[4361] = 256'h86f55afaa0fdf0feca03730740036cfb43f5d5ef8fefdcf4e0f715f94bfad9fa;
// music[4362] = 256'h85fa05fafefa2cfb6afdb300b701160144fa53f554efd8dd71d5c4defbf14fff;
// music[4363] = 256'h58f266e0b5dcbadd1ddcc1d853e64af938f75af340f813fd2700ccfca2f447f0;
// music[4364] = 256'h9ef52bfd680090017500690082fe68fed50155fbfcf7f600c60bce10580870ff;
// music[4365] = 256'h8af870f6c905eb0416f6b8f95af766edc9ef91f6fcf920f674fe6c166d1af407;
// music[4366] = 256'h26f24ded9907ce1f221ea216ae124e0ec90b330daa0fc8122a15921576188a16;
// music[4367] = 256'h3a10cc0977fcc0f80eff3cfcc3faf9fce3fb8ef89df542f76df0d4de42d8d8e8;
// music[4368] = 256'hda031d0ca001c6002709bd00e5e943e238ead5ef8ef146f00ae806e2e2f4e310;
// music[4369] = 256'h59155e10700b850164fd7d0044086a0fe80ff40f5e11a7100f0d3d0956084d0a;
// music[4370] = 256'h480b2609de0ae013921d1914c8f280e008e81aeacde8c4f6fa0b1415b20cbbfa;
// music[4371] = 256'h0bf1aefd15104013280b6507ca09dcffd3ec33eafcfff218931b1a137e0bef00;
// music[4372] = 256'h97002d09ed11501932193118f817ab1d9f2f99378233d5327636223f05391d1f;
// music[4373] = 256'h4a13101f9d352a4263361c2b4c27401a3a1052109014991a801e242c30417040;
// music[4374] = 256'h322bbd18a1126b136c08f2001511dc121a078e0f8816b317af1cfb1b271cee18;
// music[4375] = 256'h5d16bc1b56189313ac0e1c03fa009cf87ce0cdd419d8adddc5dfa9dd2bda34d6;
// music[4376] = 256'h07e041f352f952fbf904600ec1066ff3e5eceae83ae2bce618f7d80dcd109000;
// music[4377] = 256'hc3f5fcf8a30e541c6f1ec627c129a62831276225552cae2ee32d0e2bc2260d2b;
// music[4378] = 256'h3329ce1cc4174723a33197342f37bc3e344111301e153b0d3d1bcd33f741ae38;
// music[4379] = 256'h3c258816e51f393bbc48a23ba8208116a1243e320f366737af31f92b713e5756;
// music[4380] = 256'h915e6e64df634b5ba552a6504b5728591458ca4d8733a026312eec31bb2ec539;
// music[4381] = 256'h5a4ee1544a49cb2d891929182013210cc6079b08a4147c1e9c1ee215da0c5306;
// music[4382] = 256'he90369198f3371368930502a5220740f6affbc05871f30310d31682e0d2ed72a;
// music[4383] = 256'h4529ab295322e50ece01c20bb523cb345b29c30addf8a7fae60137021809511a;
// music[4384] = 256'hc71d331bb31e781f85202c2327266a260f253f23621208ff0dfea80afb1cec1c;
// music[4385] = 256'h5d08cbfd1401790530ffd7f9d608bb17621865152918d719830d8d054202d9f4;
// music[4386] = 256'h9bedb6ef43f7b2f7c2f8791a4b331c29ee1a260eb314c826c92ae92cca2d4930;
// music[4387] = 256'hcc323d32e831531e7408f007c3096b076c07040e1312e914c122182adf223a0b;
// music[4388] = 256'he7ea11eb21072b19b4160b00bee755e6cbf80c0a410d950bdd0ca003baf015e9;
// music[4389] = 256'h7deb5cec1eed65ee8cebfee81ff96a126715a30bae0e02145a0675f4ccfd1c1a;
// music[4390] = 256'h822a012548170e14dd15790a7afcf0f980f896f85bfcf5faa7f9acf854f6c6f4;
// music[4391] = 256'h1cf345f6fef7e9ffe618d227dc1ee20878fa2f04d5139e17ed147317c81b1b10;
// music[4392] = 256'hd6fbf6f6de082f1f8121200fa1fa09f81bfe22fabcf9850a7b1ee61be1069bff;
// music[4393] = 256'h7e0d8f242e35993a4e3ec73e123e9d3c0f35bb2ef22fb8392239f1244d18b714;
// music[4394] = 256'hb40e4d0f4f17001dce19cd1d05321740ed37f117b8faf8f653f879f760f7cef3;
// music[4395] = 256'h4cf69f01f00f460f88f629e000dabfdb43e0dde701f156ef54edddfc8c0acb0c;
// music[4396] = 256'h830e680e390c2a08f0048f00d6ee59e18feabef84efe9600f809ec0d07f937e0;
// music[4397] = 256'haed696d331cd1cca35dc41f5a3faf7f66bfc02fff1eb9dd765d819def0da77d8;
// music[4398] = 256'h85e42bf592faa5feb500b6f1b2d58cc3a3cda0e444ed90e9a0ecd4f5eeede0d2;
// music[4399] = 256'hc9c237c7cdc73ec094c449d569e833f3f4e6e1d4ccd99feb09f359e6d3ceb2c7;
// music[4400] = 256'h7ad84eec5feedadcd2cae6c816d7a6e921f01de478d0f8c83ad67de757e555d5;
// music[4401] = 256'hdac7bebec4b9e5b0b2ade9c197d386cfbebfa4b3f7b863c694d2a0d37ec6e1be;
// music[4402] = 256'h74b70aaacba548abb4b2a8b407b129af7eb3a3b73ab4bdb095b163b67cbb60b9;
// music[4403] = 256'h15b763b880bb8cbf96bdbeb80fb7ebb907bd10b70db753ca37dbc1d437bf61b7;
// music[4404] = 256'h04bf89c2c2c6a9cad8c858c423bde1ba4fbb6dc790dee1e353e212e3d1e2e4e5;
// music[4405] = 256'h61e11de197e9bdef4df3cbee38e7e0df2ce300eddcef2ff3c6ed30edacfc1305;
// music[4406] = 256'hd308770a890fff09a7ee01e07ee117e400e59ced98033b0aaf030504950be811;
// music[4407] = 256'he8116c105fff75e9a8e7dff8b012140e71f34aee4df67f015807b50099f6b5ee;
// music[4408] = 256'h13f2fefa74fd0000f002ef00c2ffdbfdbff9f5f9f4fb9a0153fcebe208d50be1;
// music[4409] = 256'h38fa2507bef894df0acf3adc53f9f005b4023efcbffb9af3c2e2d1dd36de0ddd;
// music[4410] = 256'h49da0ae2dcf443fc6afde0fd50fbeefcb000b8039600f7f980f7fcf8a1fb61fd;
// music[4411] = 256'ha2fe0cff08ff65fad9fb2509b302d5f135ed35e53ce10ee72beed3f356f201ed;
// music[4412] = 256'h34e350e5b4fe4e0db00cc50d6108f20785176d256621af0d60fff2053115ca1a;
// music[4413] = 256'hc91da126ca29dc26eb21e11de41abf144e16101fec26f32525196c16740df7f3;
// music[4414] = 256'h5ce981ef8a020911110a2100dbfcef02c809000b8afff6e55de071ea53ec8deb;
// music[4415] = 256'hb5e503e411ebbfedbce733df22dfdfe187e2a4f0bc069f0b0b07240504fe96fb;
// music[4416] = 256'h4701af07fc0bb306abfd00fbbc04a00a5af6c3de97d8afd305c973cfdce74ff4;
// music[4417] = 256'he1f61dfb1dfea2f650ddc4c822cfb0e529f22df08aefb8f2daf831faa9f67ef1;
// music[4418] = 256'hdbeafded7fe9dbd882d820e69df01beef5eecef75ef5b9f71105c30bf20ed513;
// music[4419] = 256'h3e136e0116ec06eeb402b20ec9033fefabe92ef83b0c021367ff74e647e443ec;
// music[4420] = 256'h8feebbeb4af3c108af106303aff66bfabf009702ad07aef80be066d978d8bcd5;
// music[4421] = 256'h2ed66ae686f851fa37fb3bfc2100260304025b003aec17db49de0cde96dcdbdc;
// music[4422] = 256'h67d96bd65eda43e212e2bce043e302e1f1e55cf86bfed8f1fee0c6d7e2e626fc;
// music[4423] = 256'h56ff12fa39f7c0faa2f382e146dd36eb2501660571f1f7dad3d24fe269f6d3fc;
// music[4424] = 256'h1bfa96f7dcf334e7acdbfddc03eb0ff6aaf73bfd80fc46f619f633fd60057d03;
// music[4425] = 256'h7d01fdf461e43bee8bf554f1d8f08df40bfc32fba50139134e140704e6f321f3;
// music[4426] = 256'h4ef689f23bef51ee81eefdeeb2f227f469f6d3052f16781571faa2dd52dd5ce3;
// music[4427] = 256'h02dda4dee9f1d0009f007dffa200d6fd62f6a6f40bf6bcea0be280ebfffa8f01;
// music[4428] = 256'h8efc66fe1807b7fbd4e29cdad7e22ae3a5da2ae662ff9f06ee02ccffb4fc2cfd;
// music[4429] = 256'h31014803d0f27fdeb4dcfcdc63db8fdfbcee3ffe8bfa4dee17e1dce01cf388fa;
// music[4430] = 256'h8ef763faab04de0335ec2dda87d73ed9e5dc40e63afd1a0b33fea7e73fdd4ee7;
// music[4431] = 256'hd5f5cafca7f994edeae9edf077f8d5f907f71b061a1c911571031304fa10171b;
// music[4432] = 256'h5916c40389fb8a01ceff74f863f751fbb9fd33017113a721061b3d0c05fe5209;
// music[4433] = 256'h51238c2b4b25250b7ef8c1fce0fad3fa0dfd69fcf1fdedfdbf0087fb70f496f4;
// music[4434] = 256'hd7f9cd0fa525ff220308f7eea7f09afaa9fd75fa7cf7d0f732fd8d11da218621;
// music[4435] = 256'hdd1c1c1a0216b200b9eefaf2dbfb84035d02c9fa85f39ef330fe20fee7036515;
// music[4436] = 256'h48172819f71d501b89138c0829078209330c470f170248f34ff597faa6f478ef;
// music[4437] = 256'h65fdd10f6812760d98123917fd0624f7c4fc300d9a1ac6162a042ff9bdff2812;
// music[4438] = 256'hc42b6c4019478348a0452e3f6338542c311f3918c322cf3367344d31a633f533;
// music[4439] = 256'h9d316935923f3a382a1e8209bb12c02b442f1622400a2afcd80cfd1ab2186804;
// music[4440] = 256'h15ef5df0d6f36af3a9ecd9e27fe119e2f7e5a2e17ae3bbf54af96ff722fddd02;
// music[4441] = 256'h33fdf9e9c1e14be3f6e170e2a1ee5e04a80fba129b14ea12ff04c5f3b6f6aefa;
// music[4442] = 256'h94f942fc88f98ffde7020907940cea0867051d0197080b2623354130ab2d5730;
// music[4443] = 256'h4331dc2f8530b029a2180011181d3332ca3e6735fb1caf117c1f32377940fe31;
// music[4444] = 256'haa1ed61a3628cb37c83a4a2df01ac425f04a00608f61655d2e551e50c950f154;
// music[4445] = 256'h52557b51cf53c852f541b32f56310b45825415571255f853054aea327527aa2c;
// music[4446] = 256'h332de525a81fb51fc71abd13ee17c31bab1d361e8c17d8110d110117561d501e;
// music[4447] = 256'hc31b5d15cc0db60f0027dd399933e52a00273b28c62a1c2d222dd61a2e0ec812;
// music[4448] = 256'h6012e80d720f322379337027c70fbcfb34ffe017d928002e8f2d5328491f4018;
// music[4449] = 256'hee18a01ee321941f2b1e0c1fea225727a3261a20c3149f13af19d40d4efa29f9;
// music[4450] = 256'hc20b461dad1f3d1bc21892110000bdf456fd3b0fd01d841a5f0121f35f05a617;
// music[4451] = 256'h9a163011520bbc088f148d29b42f8728b3285e288a2b0432fc2db42a8728eb28;
// music[4452] = 256'h472ea02d142a7325c1260628051d440d07ffeff8c8f1e3eb54fbfc0f4613d500;
// music[4453] = 256'h58f023f30bf833fbfbfb2ef630ee13f3640ae015be13d31698185710f9f9deeb;
// music[4454] = 256'hb7f89f0e48168110b6107c10a30ee515a316b217e5205523841f581e9520f515;
// music[4455] = 256'h750298000b0ed51d51200210bb0142fe1d007e005d03a813ff1fcd1e85206e25;
// music[4456] = 256'h12217f0ddefc32028411921b74157606c401a002fd01c0ffab07231a881dfa1f;
// music[4457] = 256'h7d2aed2a9e2aef26b524a030283b403e6333ca22be1cd0168514e318871ec221;
// music[4458] = 256'h951ea5240d307432bc2c512054203a2fd33c8439bd214e14df16c01d561f160d;
// music[4459] = 256'ha2ff8dfc43003416b31f1a17e40c2306eb1117246729e323c220ff1fe619d11c;
// music[4460] = 256'h671abb04b1f07fe9c5f37b0179052308c50f0b149afe28e5f8e1cde665f009f3;
// music[4461] = 256'h7ae986e1e6e10ce9e9e580e66ef8b8004ffc23fd6207440124e851dd99d8d1d2;
// music[4462] = 256'h26d516d76ed652d278da83ed12f2e1ee10f1d9f56fecc7d700d29ad3a6d288d4;
// music[4463] = 256'hf5dfd9ef95ec4cddb2d076d0c4e26bebc3e826e979e433e779f98d08990031e8;
// music[4464] = 256'hd4d6ddd744ea95fa80f73ee446d1fcd24edeabe3e4e959f21bf6fae7ecce10c9;
// music[4465] = 256'hc8d86de716e762db5cd0e1c722c044c321c74eb9c1ae50b10bb354b24daf5faf;
// music[4466] = 256'hedad9fb0f2c512d2d5cc70cc71d1d3cf50be51af72ad73ab8dac91afc8af3bad;
// music[4467] = 256'h80ac5bb150b305bcdad13adec2d02ab837b057b091ac98ac67afdbb8d1bca7b6;
// music[4468] = 256'h32b4b9b0a1b39bb5bbb10dc2f8d4f0d843dae1dc69ddd7cbadb872bf40d35edf;
// music[4469] = 256'h84d5fec14eb944c021d31cde31df91dd32dc45e0f7e4c5e864dc93c510c3efc9;
// music[4470] = 256'h55cbb3c7add583f8bb0276fc6efc4ef989fb9800760468047100b8fc10ed32df;
// music[4471] = 256'h14e812fd1c111315cb027fef2be852e46ce591e75de9d6f012ece7da40cec2cf;
// music[4472] = 256'h87e366f234f5b5f864fb3af52fe426db8ce4d3f7090072f0fedafcd1ebe244fa;
// music[4473] = 256'hd8fcb4fa39f9daf7ecf380f265f963ec28db5bde54e30de68fe28ddc0bd761d8;
// music[4474] = 256'h06eaf7f3f0f2a3f4cef565f6cff4f2f68ef326e097d34edff9f740040bf826e4;
// music[4475] = 256'h16dea3e05fde3cdd79dd64db12d904d9f7dae4db1beb1902000550fd8ffaa4f9;
// music[4476] = 256'haded05deafe12bef95ff370ab508da0d830b4f00b704f70e5d1a2e22fe1ec11d;
// music[4477] = 256'h902273219f16571191101908c100e0ff9f011903e90f0126a72943231b24142a;
// music[4478] = 256'hab2c7e284029db13a8e917e3d2f6fd08770ecffd1ff072f2a9f5d1efc7ed3efe;
// music[4479] = 256'h470f200fb3fddcebf1e7ece721e7cced72ff0e0c0f0598f42fe989f4e00c9911;
// music[4480] = 256'hbc07e80387080406f9ef49debee70efab100e5012f08660af4f7b8e29ee2abe6;
// music[4481] = 256'h4be58ce55be6bee797eb16f9ae0537ffa1ee41e837ef61e782d22ad1fbe10ef6;
// music[4482] = 256'h77f800e6a7d77fd234d4c7d909e170e5d9de23dcb9eafdfb2af7e1e26ddae4d9;
// music[4483] = 256'hd5ddd8ea2bfff116411c1a0ad8f570f12f00910e5b10f50e3c1530176e033df1;
// music[4484] = 256'h4ff579fbe5f619f56600170f95105b003cf20bf404ef97dff8e1f5f21dfc5afd;
// music[4485] = 256'hbb00b3031afa4be822e2ffe5f9e1d3dbb2e48cf6a1fd85f321e77ae412e4c2df;
// music[4486] = 256'h60db90db1cdcf9dcaaee3d05ee0360f09ddd01dcd9ec83fea700dfecdcd95dd9;
// music[4487] = 256'h4fdc79d918d9d2e655f83bfa55ed34dec8e1d9f44efe08f6b0e216db75e9b7fe;
// music[4488] = 256'hc708eafaa6e439db54dccfdc49db93e7c7f9bffc71fae4ffdf0479f795e1c5db;
// music[4489] = 256'hbadd54e16fe63de4a9e1c7df64dca4e2cdf6cb0f411e9919ad069ff9eafaadf9;
// music[4490] = 256'h6ff6faf5abf5a1fa07fe7bfec1fc11f76df6e2f654faf2fd4af9360200170921;
// music[4491] = 256'h9116b0f61ce583f61e0b980a24f815e44fe306f968081c07bf05fd0278007d01;
// music[4492] = 256'h12058b0898fca1ee4feb84e60ee391e937fd3906a2fd9ffd0cfee8fec3052407;
// music[4493] = 256'h52090506f2ffc6fe3dff43068dfe44e985e1eddc2cdc74e3a6e602e92be909e7;
// music[4494] = 256'h95e54edfaadedbe0d1e086f00801c002c401dbff83fe02f399e4a8e996f615fd;
// music[4495] = 256'h70f544e992e6aaeb84fc9f03d5fc47fce3ff6609ce0df908fe0075f9bd067511;
// music[4496] = 256'h6c039bfb610757150719ca1c8920b81cdb18011651160115e714791db018a007;
// music[4497] = 256'ha502ee0c4b1ca31e700ecdfeb8fc0cfeb5f447e7ade45ae685e830edadeb34fb;
// music[4498] = 256'h5815fb153412cd13de15e217ca115413010e74ff1efc5bf9dbf6abf6d1045119;
// music[4499] = 256'hb417a011b70dec0fbc18eb1adb17bdff71e9d6eef3f43bf8b0f7d0f1bdec5ef2;
// music[4500] = 256'h6d0df1195a0a1d03810a5c102b138916e80e70fca9f3f0fba10bf1125912c413;
// music[4501] = 256'hfe141d0e39fc6cee88f30c028f07f7fd21f14af074fe790b570aec08310f3410;
// music[4502] = 256'h9a0474f5cafab50fcf15fd1bde2bc12f3e2c2d1d180bcd146a2abf349b340536;
// music[4503] = 256'h9340cb3f3a2dc2204026c6271b1d332204386d437836951e57155e1834183c0f;
// music[4504] = 256'h230b5b1456111900a0f88dfa1d08e022fa2c1d192d05ad02f405f100e4fb2a07;
// music[4505] = 256'h08161315ab0398f2dceef1ea8be392e411f3b0041b03b4f1f5e43de847fbd808;
// music[4506] = 256'hf10299f41fed6eee4eef7ff0260049162e1b8c148912a4143316801aaf22f61a;
// music[4507] = 256'h9b0a4b080b08bb06c30c9e1c372f3d2e6e1a700b1b11711bfd1b91213e2dca39;
// music[4508] = 256'h4939b524eb1b2224bc2a622cab27de1d8c1466198923e023d033ce50c2570d4e;
// music[4509] = 256'ha940fb364d42bb53b857ba57345af45c3252163d24394348bd5c9d63c3526940;
// music[4510] = 256'h11393b369a35d73a394d975c854c122f00246a23ef20931aca1dc7330e3f4c3c;
// music[4511] = 256'hf73e0f43d441df39ba36dc2fc81bc213a2152218e01c111da21ada15d51af72d;
// music[4512] = 256'h0133b12291141f16bc194c152b0fa00bb50a9a0e9c1bbc280b262a151508d609;
// music[4513] = 256'ha60c0a0956096d162627fe21ad0926f977027f1d282a74253920341e3f17a803;
// music[4514] = 256'h58fc7a0ea522402a4823461d7c1e2c1308034e02770571fd4df78b07821e8a21;
// music[4515] = 256'h011c55191a165916211560128711d00cd30e8b21c733f430851fdd125011b914;
// music[4516] = 256'hbc13a8137215d3129a1807280a312827ed13b00f54138c13c410960b4f130f1c;
// music[4517] = 256'hf50fd1fe76fa4104b0118e13dd09ecfd4df95c03c412f713fd0459f7ddfa7f0c;
// music[4518] = 256'hea1adb15b000bbf045f19df923fb99fe6710c919ec119a0bf90ec30e6cfeebf1;
// music[4519] = 256'hd1ef9eea78eb6ef9ef0f611a020fa9fe1ef5dcf8e5fdd0fb44fcc5fbe8fd6003;
// music[4520] = 256'h0f066205d2003801c505c4078d0744050a08ea0b4e09d104980163056f153525;
// music[4521] = 256'haf23eb121b0440086a1de42bcf25301379057a0c7f29bd3f2d39502c66278e23;
// music[4522] = 256'ha01c06142221063b53407b3e80420343a340883e5c3e4d3f863dc63a0a3c8741;
// music[4523] = 256'hbf46fb44aa412c3e522f8b277724580e6d026d072c07eb09800cfe0b080c4708;
// music[4524] = 256'hd105a305f40437072d0c790eed0b6907af06e0119f1dcc19550c600044044f0e;
// music[4525] = 256'h0607f9043b10c90fb20a5008df08940e300d9f0683fe21fa9e0047051a087e03;
// music[4526] = 256'ha6f065e5bce981f8f4ff0dfafaf924fcc3fd3efe44fcd4fe53fb94f96cfa4af5;
// music[4527] = 256'h70f676ea8bd5ddd549dab8d850d9b9dd5cde75d7f0e176f62cf68af300fc4e01;
// music[4528] = 256'hbc05380bb909ff020a05e80b66061401aefbd8e829ddc7dd6be0bce08be319f6;
// music[4529] = 256'h860189fd3cfb7af592f51efc9efff7fdd1f40bf560ec83c8b5b535c1c0d0b0d7;
// music[4530] = 256'h10d789dbf4e09bd310b865ab8abcfbd34ddc6bd9a7ce88c5c0c6deccdbd2fed0;
// music[4531] = 256'h07cf80cc09b982aa51b0cfc0cad232d103c01bb0f9b01ec6f5cefec905cc70d0;
// music[4532] = 256'h54d3dcd1b7cde0c173ae6aa94db0f3b2d0b5e4c162d4e0d88cc866b726b1eeb3;
// music[4533] = 256'hdbb68db838c8ddd7f0d6add725db16dbcada14dd13e087d149c173c263c186bf;
// music[4534] = 256'h91c1dcc39dc5f1c044be2dbe09c5c8e0edfcb70002f684f323f2f4e3dfdc06e7;
// music[4535] = 256'hc9f7e2014cf623e62de722eb4de507df63e90e007a094000e8ee16e608f19402;
// music[4536] = 256'h6e0e9b0a2dfa57ee83debdcd10d2d2e31df045f317f48ef5e5f59af5c6f56fef;
// music[4537] = 256'h75da88ce97dd3ef3f8fa1aecb9d613d185d5a1d8cbd619d6d7d59dd41ddf3def;
// music[4538] = 256'h40f3dbe723d99dd539d53ad189d2b8d86edae7d8dee3edf5c0f349e1bbd4afd1;
// music[4539] = 256'hbad2add470df49f33efab9f184ed75f3fff2dbe3cadba4dec3dbabd965de4ae1;
// music[4540] = 256'h6fdf9ce7a9fb3c03d0fff0ff2efe63f3abe2f7dce2ddf7d660d89fe9f702df18;
// music[4541] = 256'hc11c6619e3138407920317056101410186094f1a1c26141e440d8f03bf0a531e;
// music[4542] = 256'h3c2b8329ce1a940de214582420282925801cb90fa106a9f970ef4ef55702de0b;
// music[4543] = 256'hf6053ef555ee00f9410e5315c305b5f25feef9fe530f380c30f9bce6dbe82dfa;
// music[4544] = 256'hba0bb40e38fb8deaf3e9ceeb10ecefe95fe779e997ee49f209ef4ceac5ea11ea;
// music[4545] = 256'h69f27605690a92fecdee01e708e681e3fbe837ee7ee8c0e0e8db31df53e5dfe7;
// music[4546] = 256'h64e8d6e835ec75ee2def87ea16e566e511e89dec89e43ada09dddee21df5d800;
// music[4547] = 256'h21fceef77af2bff51af9fcfe4b0f9012ca12ca09e8f3e9ee4af47cf732f651fd;
// music[4548] = 256'he811d51788152a181315d310b611af152019b91ad71b0a1ced170d14aa13ac07;
// music[4549] = 256'h4af8dffbbd0576070b0318fe63f934ec18df34e552f94c06d002fafa64f9aff8;
// music[4550] = 256'h72f8b3fa0ff51ae659de7ee8c5f974fd56f0bee177de76ebe5fc6bffcbfaf3fa;
// music[4551] = 256'h8afa25fc49fc7af578f159f2e6f7ecfd90fe68fe5df80cf256f3edf34bf912f6;
// music[4552] = 256'hacdf5bd4f2d6e4d69ad4afd642e648f54ef75af8e3fcbbf81ae5a1d75dd84ad8;
// music[4553] = 256'h25da3ddcacdfcce449e46ce3e7dde8df20ef1bf58afb1f026e05b60ee50a6c05;
// music[4554] = 256'h150e3a13b712400efa0c45149f183f1aea17330627f030f08d04c21489118a05;
// music[4555] = 256'hcf027007ea12ef18810cdeff64ef2ce6b4f608fef0f989fdd2fe28fc87f9b0fb;
// music[4556] = 256'h8ef6b6e5c3de01e758f609ff3400a0ff80fafcf858f9ddfa8afe16fcc2f90bf5;
// music[4557] = 256'ha9f3d4f803f048e562e4d3e047dfd8dd19d87bd74cda40dcc3dd91d957d70fdc;
// music[4558] = 256'h41e139e290da6eded6f2abf939f531f5fcf746f0eedee4d993deb2dd19da1de6;
// music[4559] = 256'h9ffacbfce6fc6300b8fdd8fa4af567f30ff475f88afc1cf0b5e3cae5d3f541fd;
// music[4560] = 256'h90f5c5f828fb54030e1329122812ca15151819199817d81ceb15e10259f875fc;
// music[4561] = 256'h7b0b0514490f5902f0fb1f05ec13f41cd4153d07d6fed80a501c1f1199009500;
// music[4562] = 256'h5f0415081c0cc10b9ff627e23be5f9ec02efceeea8f9a4055600e9fe9f092e11;
// music[4563] = 256'h920d2a0d56148017001bf6100cf81deef1f1b4f469f421f334f156f27ef61df9;
// music[4564] = 256'hd3f94ef758f4e2ef7fef76f4b0f6880588131510cd0cdd0a4d0a2801c7f3c1f5;
// music[4565] = 256'h52fd4c09260c04fce1f1f3f8b30de01bf31ae1169c12de115e141d16bc0cd3f6;
// music[4566] = 256'h35eb25f419077c1083111c13060fee0ea911d20d8e14342378283629a8289823;
// music[4567] = 256'h641d2016b616ff24d931a330592068125e1324173a1a501da820b822d323e728;
// music[4568] = 256'hc229fa2c1b3f934d773f21264326d123820f270a140bd5094009df0f70236d2a;
// music[4569] = 256'he9238518dd110b17c614b918fb20e62108273d1a4507670204fa8af4dcf2adf1;
// music[4570] = 256'h82ed4ae9d1f690029b00b3ff61feb0fa30f6f3f9effc90ed2fe04be6c7f87b06;
// music[4571] = 256'h4c008cf052e9b3f11d031e0c3a0563f691f1fd01e4153c1baa1dab229722231f;
// music[4572] = 256'h201ea5230321a011dd0f1b1d8c29732de62c413504369623c213201647290035;
// music[4573] = 256'h5d33a13f46545652bb3bfd2d0131e73546388f372c3603399d3b8b3bc4399337;
// music[4574] = 256'hdb355f36c73b563a2334f13e5a537c5b2456ff549655163df420e71c2e1de61a;
// music[4575] = 256'h3d1da3293a3a5f3ae52d7a23e9202e1d4111f81263296f3a6833081ee40d0c11;
// music[4576] = 256'hd7268a329931c633ac30522d112b7e283d2b0a2b572cd42e652fa8311d267e0f;
// music[4577] = 256'h3105990d211e9626881d930c48077b118c20cf239f16130bf7077e052c00fc03;
// music[4578] = 256'hed18ee2b5028a310bbff8aff1201eb01b1022f07c608cb0a2519631caf176819;
// music[4579] = 256'h70170319711da5247926d31f381c670e1709ca163c19f117b7187b1732192b1b;
// music[4580] = 256'h7e1bb61696131216d4169117d820d12f5e305a22ba170d179c1936169a19672b;
// music[4581] = 256'h9f3c5e3bf325561735143a0860fcb6025314931d531dba1db61d44183313c612;
// music[4582] = 256'hd90b98fdedf63effb70c1f125a155016e71262116712f8158f12320c6a086afb;
// music[4583] = 256'hd2f32df782f9bdf790f58000da0eae0fe3048af737f697003e0db70d8a0046f7;
// music[4584] = 256'h23f636f5b5f0f5f88a0c5514f8148f14491ada1c000c0c023005e3045803e10b;
// music[4585] = 256'hf81cf4211b2265254425d527a7289f26af1a6b0b850f251c6527cd21a10a6c0d;
// music[4586] = 256'he222492b702d7d29411ea1176d1a1322e424602963383a40043710253c189221;
// music[4587] = 256'hb035a040f4390b24a81ace28443a284159344e155b032b11e820852211200921;
// music[4588] = 256'h9a24fd1823093109930d3b0fad0ceb0c2c092c02cd10bf2052221322211d6c17;
// music[4589] = 256'h5e14081a321af50348f6d3fba2ff66ff23fde6f47ff0f3f564f427f17cf086e5;
// music[4590] = 256'h9fde03e0d0e373e9cdea47e9d8e6a2effc00700261f654e816e47cee7ef7b5f9;
// music[4591] = 256'h95fb79fc67f7d2e759d6cfdb4af5a00001fd1bf958f401ee58decacd90d2f1e4;
// music[4592] = 256'h23f0a0f1d5f2e5f5cbf47ff4f3ffde0873048006c40da70db30b2e04dcfc47fb;
// music[4593] = 256'hbaf08ce730ee6bf20deafadebcdb17e0d7e448f190ff4ff8ade27cd5f6d95adc;
// music[4594] = 256'hc0ca06c234d0d7db29d5ddc065b16bb2f0ba71bb9ebf37cd2bcd62cde3d414d3;
// music[4595] = 256'h63d238cfe5ca74cc8fca4ccb37cc25cda0ce9dc1d1adc2a8c1b77cc831cdadcd;
// music[4596] = 256'h80cd8cc984ba87adebb07db208ae4db238c3efd181cab5b779ae22b07cb1b9ae;
// music[4597] = 256'h9fb541cba8d88ccc61b7afad89b982d024d6ecd1d8d24bd21bd419d929dc50d8;
// music[4598] = 256'h17d556d804cf47c022be0bbda5b706ba7fcc13e0cce0cdcd1ebebdca55e5a3f5;
// music[4599] = 256'hfbf572e796db2edd50df62dd93e254f067ff270268f4fdeaa0e94ee59cdfd5df;
// music[4600] = 256'h2fe933ed9cf6fe066a026afe710174f8d8f24ff193ede4e1fdd2c8d4f7e1def1;
// music[4601] = 256'h3dfa36f03ae335ddddd65cd2c3d622da14d8f4d7f8d898da85de21eca9f9d0f0;
// music[4602] = 256'hf0dd90d4f4d530d7e4d11bd956f032fe0efb0ef752f50beb16db7cd6ffe4ebf3;
// music[4603] = 256'h07f60ff3daf3ccf875efe0dea4da6dd94bdaadddefe2dee4f0dffae956f5c2f3;
// music[4604] = 256'h6af5d1f85afd0bfe68fbd4f4bce09fd6c3db4cdd25d8aad875ec74fcbef706e8;
// music[4605] = 256'hb1da94e19ceff2fb2805edfa7cf2b0f79bf689f3b4fb3d0c6314e70baafca3f9;
// music[4606] = 256'hbe0b291b371c211ea1237824f3193f0d790c1e18f7249627232967259e10e1fc;
// music[4607] = 256'hcbf234f5f8049f111e0eeafbbef069f2eef4eff77bf737f746f6b7f62afbc2f7;
// music[4608] = 256'h22fd170c3e0c3900a0f1c0ef02f477f043ed77eafbe9b2ec94f8da091f078df5;
// music[4609] = 256'h36e70ae4d2e5d3e363eb2bfc46099d03a7efe2e8a8ebeceba6e890e605e9cfe6;
// music[4610] = 256'h83eedaff84062d07fa068b085807b5053b0af9ffb7ece7e7d0ea22ea48e694ec;
// music[4611] = 256'hfafcdc0244020409480cdd0098eeb3e777ec96e314dbadf3c40ee40dccff34f2;
// music[4612] = 256'h46f0a7f682f6daf8c505790dea09cf07290a9607bcfbfef167f8c2062a0d380c;
// music[4613] = 256'hf00c5b0d5a0424f87aef60ed7df803fd8deb4cd9d7d7e9e84afdfb0071f38ce1;
// music[4614] = 256'h98dd88eacafa60ff1cf26ce5fbe4cbe452dc6ed773e98dffb5fddeea26daf0dc;
// music[4615] = 256'h23f049fe0ef886e391da66dd02db1cd541d947ee23fe39f62ae53adb26d966d8;
// music[4616] = 256'hc4d89bd91cd9b9db25e066e251e114dfd7dd4ddd16dfeadf1fe256e6e9e0c7dc;
// music[4617] = 256'h6eeac0fb0afc6beb63ddefdaa5db89de44e31be42ae0fcdcf8ddffdae9ddf6f2;
// music[4618] = 256'h17ff60fa1ef7a0f44cf7fcfa03f63cfb7d0d9c155815af156e137f164c19b914;
// music[4619] = 256'h2415551595147115d5166c1e9b1dd41b2d18d501daf611f4b8e797e1dde3a4f3;
// music[4620] = 256'h1b02220358023a001902e005f707e100fbea79e151e585e674e7a6ee5f01130a;
// music[4621] = 256'ha1fe18eeeae2c3ec49fe3e013800c300f3ff75fe6afb95faf5f9f7f6a2f850fe;
// music[4622] = 256'h65059e07d9f633e0d7dc91ed3b00c3ff16edf8dbdedf05f445fea6fe64003b01;
// music[4623] = 256'hc0fb06ebf3e046eaf5f7eeff3afab5ea29e2e8dfc2e068e470e7ade781e2cfe7;
// music[4624] = 256'hcaf989ff81ff310144fddefdd500ff010c091e173f1ecd0ee5fff2ffecfd35fd;
// music[4625] = 256'hb9ffddffcefd60fa36faf4f96ffe8c0df11a5c19fa0af601fbfdd3f5e6f456fc;
// music[4626] = 256'hb0027e0050f920fb84ffbdffed00a6fea0f50de928e7b0f62204290573009bfe;
// music[4627] = 256'h38015d012004f804b8f574e580e7f2f734059b06c4056805d501b3046c13a715;
// music[4628] = 256'h1a02d7f7d5fd97fee3f5caf47c04bb0f1e0f650f55102f0adcfaecf41100ed0c;
// music[4629] = 256'h9812aa0945fc04f713f408f1ebf259030315a514f210a3144015e40542f129f1;
// music[4630] = 256'h47f9b6f55bf8530be918a218f21a80234821c00c43f9c7f8ce067712ca0bd102;
// music[4631] = 256'h9d09f112051e5328fa20d011240bfa09c5076708f5108418ae18212061330a3a;
// music[4632] = 256'h412c4d1c5615b71d86304638952b541c641bd7217627af27b11d2616e41d472e;
// music[4633] = 256'h583716307c22811bb3134f07c303d1051608350c240b030a6a098407910075f0;
// music[4634] = 256'h2afce9187c1c0a1f2c24a922ac1c2808fafdc6001500bfff0df789ebf8e562e3;
// music[4635] = 256'h6be56ee881ebcdec45eab4e641e529e393e231e8a4ea1dec62ea70e832f99a06;
// music[4636] = 256'h920a4f130d15db158918441b281c0f186919a0143f07f203160e6f1de0209919;
// music[4637] = 256'hd312bb164b27c831902c4123a72d1c42db450e4664455b444b486e483f4c6c50;
// music[4638] = 256'h944d9a4a8048cb49174d60524e52b04330358d381046474b6b4d2e52f5545951;
// music[4639] = 256'h833eb131d72fbe23851f2427282b8c2cbd290c24331d8b1baf1c7219eb238b35;
// music[4640] = 256'h0d38e938513c0e3aaa3819351f31ae34c7378f371034402e7e2d8a2c332a3e28;
// music[4641] = 256'h191f9815be1523162b119817542b2933d32cc12745222c17040c0c0c2d1b3a2b;
// music[4642] = 256'hfc2c98259f22e225ee29342cb627bb18d9083005a012232185210821d6219a20;
// music[4643] = 256'h7c25a227ef2614255e1e381e9a1f001f911d570e8c021507d510d522d6282f18;
// music[4644] = 256'h6313e1208533ba3b642a0f177f12311594161312261ad82a722dbe28102a0d2b;
// music[4645] = 256'h2b1e9e0e9f09c2098f0a700d401bf21d8f105a0ef30b810de814c8118110990c;
// music[4646] = 256'h510d8b0f16ff93f707fb3afa9cfbc3f8adf4a8ef86eaaaedf0ee49efe5f34df4;
// music[4647] = 256'h7afa3d099a0d2f06aff5e4e840f4d506a00b40ff38e9abe06aedcb03100f2e07;
// music[4648] = 256'h12f87eeeecf38dfec204250b640fb70c12035bfed9fad2f0e9eb77f1cd001706;
// music[4649] = 256'h3bff3805640bf209f407d80554033d047c197b266e155c0e9713e11360128d0e;
// music[4650] = 256'h150d89101212d211921c7f2a192a7b26962632268d285d2c962929262b30ac3f;
// music[4651] = 256'h1e47b9462c47784315314e24a3251328d328be2b193b004698421e40f5350a29;
// music[4652] = 256'h9a28b32cf028311ac011531acf29d22f7d2e1b31172ea929232aa3270129212b;
// music[4653] = 256'h662ba92c5d2c7c2d112acf257627c51ed20eb70ea81ee72dc32fd21ee40be20d;
// music[4654] = 256'hf41d162815251d1bb6112a10ef19eb205b1e421d4f211c1aac03e0fa38f7b6e2;
// music[4655] = 256'hfad8eee3c6f1c1f7e0f6e9f920fbdff901fbe2f8c6f519f352f113f042f06ef2;
// music[4656] = 256'h5fe88ad823d6e8db5ee0f9e0badce8d4a2cd43c984caaed79ae485e513e683e6;
// music[4657] = 256'hcae1e1e75efba405f1fb03e88edcf4e6e1faa8025ffa8eeaf3e03fe85cf6adfc;
// music[4658] = 256'h1b01c3043effc6f6dfec7dddcad5e1dc77de70cc42b807b61ac796d921da43d3;
// music[4659] = 256'h16d22cd0f5ce5cd0e7ce9ecbf2cb6dd0c3d1bcce73c5e7b2f2a93eada4aa73a8;
// music[4660] = 256'h99a84ea6baa8a0adf6b0fab0ecadd6a64ca09aad7cc382c925c477bde4ba4bba;
// music[4661] = 256'hb1c0e5c8edbeeaaf71aa63a8eca566a8d1b8eec68ec86ac60bc492c336c380c6;
// music[4662] = 256'h67c885c77dcefccbf4ba02adb2ae12bf1ec9f9cce8d2c8d410d6c1d66bd6f1d6;
// music[4663] = 256'hf8d576d588d5ebcc86c570d431e8b6eddfec37ed62eeebe247d4cfd6aee6b0f6;
// music[4664] = 256'h06f360df11d272d8afed81f752f4fbf32ef8c8fb3efd88f975e1e1c68fc31fcc;
// music[4665] = 256'h29d02acdcdd2e8db51dfc1e73cecf8ed04e98be0d8e3e8db28cebfcf93d2a3cf;
// music[4666] = 256'h88cc2ad98dedc9ee6add58cea4cbc5c9f8c695ca45d23ed9f4db2cdcead339d0;
// music[4667] = 256'hdbdedae887e9c4eb4ded10e880d53dc794d05be503f01ae954d8d8cf38d919e6;
// music[4668] = 256'h55ea73e9d9e91aea85e086d4dcd42be309f3a5f05de005d5d9d428dad9d697d2;
// music[4669] = 256'h1ee0a1f0a7f4b2f590f22aeae5e8a5ed88f0c7ed09e7abe8fdf81f0a6e0691f3;
// music[4670] = 256'hf9ea76ed53ee12ee31f030f212f177ee57ec6aed09fa010fb015330686f3aef0;
// music[4671] = 256'hcff7fcf674f403fc0303a1044f0ecd1c301b6e0eed028d006d100a1cba17f415;
// music[4672] = 256'h2c1a3b1c961253067d036c03bb00d1fc7effc204bd0d4f1e1a215f1797117912;
// music[4673] = 256'h9317d319731a630f7efb0cf7e5fb8dfc01fdb905bb14001b98180b17db136508;
// music[4674] = 256'h90fc63fa36fdc9fd0efe51ff0dfb0cfd710f6f1cd9181607ccf4fcf6040ab518;
// music[4675] = 256'h8715cb11dc178a142405e9f4c9f7c509a10fe10e5b104311120cebfbf4f38901;
// music[4676] = 256'h8d1b1f2b9022a213e30e8f13cf1a721eb5144cf902e960f5fe03b20306ff4201;
// music[4677] = 256'he90361f991ec16eb87eb6fece4ee58ed3debcbe7fce96cf393eddbdb27d6e2dc;
// music[4678] = 256'h1ade67d6ebd8dfe674ee5ae7e5dc5de08be5fadf3bd9b2d2dece85d265d90ade;
// music[4679] = 256'h9ade23dd14d758d2dbd6bfda4bdec6e7b7efd0ee7ce4a8da1ddcf6e8a9f2aded;
// music[4680] = 256'h87ecdbf4fdf1b7e107d3a6d101d2b6cd9fd886ee74fa13f294dbcdcf54d572dd;
// music[4681] = 256'hbde0e5e751f1c5edd4ea0cf1a4f225f393f4a7f529f6d7f3e4f229f06bf0c4f3;
// music[4682] = 256'he7e91edfabdee6dc6ed9fad722dbbedb41d9d2e5ddf23aefade593d9edd812e9;
// music[4683] = 256'h8ef5f5f2cfe25dd72bd6b8d321d6a3db6bdd8de18ee580e3addee8dc26dc08de;
// music[4684] = 256'he3e461e7cae8d3ecc4eb20ecdbedb5eb5bed3bed90e675e4d5e66fe6c8e674ee;
// music[4685] = 256'h83f6e3f539ef07e5fadc4ae076ec5ff247edfce8b7e457e33febb5efcff08aef;
// music[4686] = 256'h8de9bfea04ede5ea74eafae56fe1daea9bf976fb02f65dfb0c0ae40b9703cc05;
// music[4687] = 256'hd108560b7a091b005004b00051f641fe890037049e0ae609730ed6049afa9400;
// music[4688] = 256'he8fb16f760fc4a02440d0b16c511fe05affb33fa5e02b1054d0245036802b1ff;
// music[4689] = 256'he9fed1f879f3eaf045ec88f09cfb500637124f101b0251f132e1bee6c7f277f4;
// music[4690] = 256'ha8fa0ef76ded0fecbceadef060f646ee14e8c9eaa5ed6cf27bf947f6d4f31efc;
// music[4691] = 256'h9dfff4f960f339f82b047e038ef22fe0a3e1eeea69ec79ed2cea58eb08f355f2;
// music[4692] = 256'h82eea0e793e50cf438feabf9a5fc23065a019bfdd4021d06400d780e670ddd0c;
// music[4693] = 256'h38019b08a819e11c74273921a011641d1124ab23532ba92c16311437303b1044;
// music[4694] = 256'h9b474747ca4906508c51e944e53aad3a6c3c7641c448aa502e52bb4e3e505754;
// music[4695] = 256'hd9576f518646db4d93573a5222519c56a251cf498e4cb54e51483948a1529c52;
// music[4696] = 256'h15495f4a024c2b4b8e50a44e4646cc3f02416849c54cbc50964f124acf51e550;
// music[4697] = 256'h77447645a54d9c4e3e49e248ce48f8401b3c643d2640503c7a39fb417742563c;
// music[4698] = 256'hdb3e413c1d365f39773b3a36e3310c2f862b6f2d1536ab3837371a3a6634c22c;
// music[4699] = 256'ha5302f2f1e21c81140129e22922cd92acd2643274528082409245f291c2bc123;
// music[4700] = 256'h5b19df19da22b225f51c1119a4222727aa255c27f4200e1480174223f621c520;
// music[4701] = 256'hf81e7816141ffa2c2c25d7199f113805100ab0197e23b82e75266614b80ea606;
// music[4702] = 256'hdf08400ae8046f10170f15055708e3050ffe71f064e70dee7ff284f3b4f0bde6;
// music[4703] = 256'h22e0dce3c5ec7ae809daded726d7fbd05bd95de104db38dedae139d890d582d0;
// music[4704] = 256'h3ec16bc5edd0b9cbccc860c227b4c4b591be33c611cccbc917c73ac4cdba91ae;
// music[4705] = 256'hc5aeccb665b6eab831b948b44db6fcb311b386b8afb89cb7e6b860b984b35db0;
// music[4706] = 256'h85b7dcb990b880bdebc291c2b9bcabb670b54bb634b721bc57c264c5e3c256bd;
// music[4707] = 256'he4bc90b911b4e4b453bac2c8b1d1b2cb00ca69cfa1d128c9dbbd08c1deceabd3;
// music[4708] = 256'hb1cf24d1e9cd85c8cecd56cbd3c4c9c8a7d1fed569d195d568dddad5b5d0cbd6;
// music[4709] = 256'hb3db54d8b8d53fdc28ddd7d385cf94d627e034e5cae444db75d44ad7d6d482d2;
// music[4710] = 256'h3bd850de01e8beeba0e332e44be693df2edc7cdd42e644e8d7e16de717e32bdd;
// music[4711] = 256'hf3e70ae41edb80de84e5c2ead6e5fee773ee89ea96eaf8e54ede1fe5e3e9fae3;
// music[4712] = 256'hc2e01ce4c4eb72fb73095b067bfe77fe9cff55fef0fa63f960fe7e02de038808;
// music[4713] = 256'h280a9d0a870afe03a605df0b4e0f8412600435fbdf08d90c2f092407ec05650c;
// music[4714] = 256'h1509e101cc05d706d10c5a0f1c02dc05d6119f11f414ea0cf5000d0666095b10;
// music[4715] = 256'hcf17710bc60198022f015d0b3617270af8fcfb012a07500743024a0260077108;
// music[4716] = 256'hd80e600820fec508fa0803027904c206b00a8b05b2febaff45008008810fd40b;
// music[4717] = 256'hcb065a04ff079c105416fc11ac0ac407c1026702040bea0fb9093704090a000f;
// music[4718] = 256'hf50bd8ff7ff50dfd140497075a0d080b880eb8116707abfd66fc2e00d5fd39ff;
// music[4719] = 256'hc009870c7608affd10fd9f09ef0834059905a7065a075e05ee0b920638f99bff;
// music[4720] = 256'h180246fbaefba705790e92073204310abc075101f2ff2603b6fcf9ebbae463e7;
// music[4721] = 256'hc8ea6bee9cf070ee86eb4aed8af1d5f701fbd0ef1be454ea86f170f157f3d4f1;
// music[4722] = 256'hc4ec9ce495ddb5de9ae05bea62f04ae48ee320ebcfe5cde516f367fcf2fa6df9;
// music[4723] = 256'h28f759f235f6d4fe0f03f80926154c15240db008e0fe06f809fd6d01af054702;
// music[4724] = 256'h6af474f3a1fab7f68ef7e0ffbef9d7ef9ef2a5fc370314fe8bf953fc74013506;
// music[4725] = 256'hfd060711c11ce31e5527d627a521d424ae23bd2d9c3bf02d19250a2aa1274331;
// music[4726] = 256'h013ad1307337f1448a405e401a4052360e3ba342193de73d234228434346f63c;
// music[4727] = 256'hc32f2634673e3949b7518b4d2c497445ff3b353c41440b474f45c841d13fa040;
// music[4728] = 256'h59408340a9454746143de5321d2b962c942cac24092a612e972b432b5f239d26;
// music[4729] = 256'h0029bb1ee0280e2d3320812338296b2827293225d11e101d871f0824d626e722;
// music[4730] = 256'h7c21a321731bd01b921cab18af1baf1ca519bf14f7134f1ccf1a271a69237f23;
// music[4731] = 256'h532404249a1a671671149714a11581129b187522c121cb1be512940c0210300e;
// music[4732] = 256'h2c07220ddc129710cc0ffd0cfb0f0519851aa6126f0b980eff0e03082b06d606;
// music[4733] = 256'had0a9a150221f31d72114d0c980783033c068b0ed0172f16780f8405c5003b08;
// music[4734] = 256'hf2078d0afd0cf302bf097f13850f7f10b8081df747f7e3025200aef7d3fb9b01;
// music[4735] = 256'h7e02f4044703cf030107b3f8cdebd0f3d4f870f9a6ff9b03e7fcc2eb8be145e1;
// music[4736] = 256'hc2e34fea12f04ff226ecd7e51fe5cedd5fd930d81ad659dbb9d9ead7b1d9d9d1;
// music[4737] = 256'he5da75e85edea6df35ea39e848e486da07d5e5d913db55dc2ee087e1abda4ade;
// music[4738] = 256'h39f367fabcfe2307b0fcc6ed43e620e480e701eea4f2c5f318f5c6f0a1ee3df5;
// music[4739] = 256'hfbfac9faa6ed02eaf2f1c4eecbf334fabeeee8e70bee92f105f5f3ff5efd50f7;
// music[4740] = 256'hf8fb5ff7cbf948fedef65cf8eff89af96affa3fbfdf457f1e8f48cfe0905a803;
// music[4741] = 256'h28fdf5f773ecd6e1b2e2e2e0a0dbd3d781da96e477e7cae2d3e10ae892ee93ee;
// music[4742] = 256'hdce9c1e39ce78def71ee22f42ff3c3da41d3ebdf8be27fe132de79d9e3d6c6d1;
// music[4743] = 256'h99d2c5d080cd7ddb8fe86ceb05ecb1e3e1db91dad2d767d7bcd7c8d9abe379e6;
// music[4744] = 256'h8de441e81ee44ce340e7fedf0cde5ce01fe2f1e578e294e5b4e559dd13e8c6ef;
// music[4745] = 256'hb6eab1ed7bea71e6a9ed69f27df21eecf6e3ffe51ee8b1e9baef15eb6de448ec;
// music[4746] = 256'h94f183ea8ee246e3cceb47f2b4f659fa97f662f10ff056ee8bed10ef11f056ec;
// music[4747] = 256'he4e97cf2acf771f296f3a4f4dfeeb8f276f547ed8beef6ef27ed1bfa24fe59f2;
// music[4748] = 256'hfcf1f6f43ff7bdf12be0d7e27af180f600ffa0ffe3f268ec78ec0cf191f70ef5;
// music[4749] = 256'hd6ed39e8fce619ee05f054f0cffcf5fd2af1d5ecf3ef35f97efd94f654f44df4;
// music[4750] = 256'h0ef1a4eb42eb15f6faf62ff318f844f3e3edd2ee35ea84e35ae64b00b6101608;
// music[4751] = 256'hc10cec0ee50415023bfc16018f0c350a4b0a720a0d065405df04580b6b11b80a;
// music[4752] = 256'h460a1d0f4b0773ffe7fda6fe7e03f10979137611eb04900427068906d209e50a;
// music[4753] = 256'hf20e4e0d640b3a115d14c70fc0fe25f85c02dd037607a90cf809480c710fb80a;
// music[4754] = 256'hf0fcd2f0d6f062f359ef44e709e70be8a9e225e507e619e1b2e163e36ee912ed;
// music[4755] = 256'hc0e88dea4cec7cec71f33cf241e894e99df482ffde03cd01230564075f04470a;
// music[4756] = 256'h6e11030aa6fa83fb9c05caff9af794f5b5f8cefe82faaaf95efe90fc9df546ed;
// music[4757] = 256'h0ef3edfaeafdfe0afa0d07032afd8cfca70040065209d30b2f0c5d09a90c1415;
// music[4758] = 256'h521b481a6e10db15b123231fd41d91208e1a7a19e723e2341e3b47399642ad4c;
// music[4759] = 256'h404b43452c444145b5421843a049104842449a4d94530753ac4d6b400744b84c;
// music[4760] = 256'h514d1b574f5b2755a350a84aea47f94a114a9348c44dd04e735366573a4b8f46;
// music[4761] = 256'h104759449c47f547b94bfe4d3c46e94096427c45b0447a4bec4e134b924c4c41;
// music[4762] = 256'h363bc5415e3c963e3b467446f5466148614b9544d934112e9833233bef391e3c;
// music[4763] = 256'hd347334aae3dfe2e772685287d31ad355b349a350a409e4a97482f4af14e7549;
// music[4764] = 256'h5547014494372335a0391132cc257b23182b9a32a52f952d682f3b29d2259a25;
// music[4765] = 256'he3210820c51d6e218d2567228026e9283020531bb41db424df25bf217427bb25;
// music[4766] = 256'h8b1ce41cd6164216d5200523b9201f167212d11b40158b0e6014d810920091f4;
// music[4767] = 256'h89f6fbf7fff0e9e9eceefcf997f640f4fdf6acf0f7ed1deb9ee759ec8cef0ff1;
// music[4768] = 256'h09ed88e3fce11de693e82ee3f8de42e2fbd96ad38cd9ddd334ccbed15cd2f9c8;
// music[4769] = 256'he6c8e4ce92ce68d608d35cc306ca1acb4ac473c375b6ddb7c6c45bc577c58dc3;
// music[4770] = 256'h8bbfe9bc66bb6bb76db73ec02bbcdeb584b809b407b4d7b6c8b254b4a7bce6bf;
// music[4771] = 256'haebe4bbdeab5e3b597c089c039c20cc802bf95b433b386b545bb57bfd2bfdfc2;
// music[4772] = 256'h52ca69cc45c72dc507c273c38ecf30cc6fc3d9c9f2cb2fcdd1ce4dc542c3a3cc;
// music[4773] = 256'h7dcf0ecf76d5bcd5dad2f9d6a1d239cc29cb32cd1bd63fd510d5b3dc94da15db;
// music[4774] = 256'hfbda52d3f8d177d5dddd53e257dbebd73bdabbde26e3e0dda7da8ddfcfe018e5;
// music[4775] = 256'h9ce672e5f3eb3ee26cd51adb11dc5ee1b5ea1ce15cdc64e8f8e988e616ed3ae6;
// music[4776] = 256'h80d997dfaae528e952eee0ebd7e7fee503ef9e00ed07b907d404a50020024704;
// music[4777] = 256'hfefe0cf97efa82fd02fe1d012c0960119d0e9c02c4ffde06d507c5061b0f6416;
// music[4778] = 256'hf212040d4406f3febd008d07300c1d0d000b980db407affd6606330cf905f001;
// music[4779] = 256'hd1016d07160a760db30d1d051d06d5087e0b4e110a0ca2010ff2e3ebdff38fec;
// music[4780] = 256'h02e40ce3c5dfabe73ff0cbf502046c0c9709a907ac0b2110770f3d09110192ff;
// music[4781] = 256'hc901be05c40c3808d7ffd70394092d0a04063005150aa60b510cfc07f6fe4dfe;
// music[4782] = 256'hb4061d0d280aa10ba81165102a0ed50ad3070001d0fb8d0510066800c108f40f;
// music[4783] = 256'h2710d60772ffff02da07740736099d0ce3080207930697022a09280a58043a03;
// music[4784] = 256'h4bfe3102f00216ffb107bb051002960469fe4bff0408b90bde0b4a0de009d903;
// music[4785] = 256'he506d50644095a0f6804be01990d930c4d07ac06ea070f0d4802b6e884e7c1ef;
// music[4786] = 256'h51ea21f113f750f5d7fbcefb71f64df124f039f143e744e65aedb0ebb0ed11ee;
// music[4787] = 256'h70e77de44ae46ce3a8e4e6e68ce6bbe5c7e719f28efa3cf63ff261eed3edccf5;
// music[4788] = 256'h70f846fa3602ec0a510e9e0ce80c190cc90e3b0e3006af06a404f5ff35febaf4;
// music[4789] = 256'h66f4c0fa61f83cf694f467f52e05be1655140514cd1bf0131d11881699164a1e;
// music[4790] = 256'h4825372a222dd124db203823d8225e25462b8f2ccb29c42eb034ab32d2348037;
// music[4791] = 256'hb7345739713ccf3ab33ffe3b75385440ea3e1a406a463742a73ee543c64a6c47;
// music[4792] = 256'h51426d42bc419244d14254442f49bd47194b1e3f382cde2996244824c0261e24;
// music[4793] = 256'he129ad2bb929892ff42d7b23c725fe2808211e22c023c924762b3427f5241928;
// music[4794] = 256'haf250e235122c3224c2210272c26c619b71b6b220f201b1f401e8a1deb203b23;
// music[4795] = 256'hdd1efe1f5427412386210927e321081d661fbb1a301cc425001f8d18511c431c;
// music[4796] = 256'h5f22bb23991cbd1a8218641bc41d0e16860f100a1f0825126b1f4c1f9714e20e;
// music[4797] = 256'hbe0d34087803dd0bbf12900f5a11ad0c4c08420f7d0afd09ed1480141e11d60e;
// music[4798] = 256'hba12a7161f09d505380f5f0f18119c0cc402e804470c5a12840fc307e103bd01;
// music[4799] = 256'h7807e10a490a800c3d0208f8b4f89bf7b5f6a1f72cffbe074a042f0088ff96fd;
// music[4800] = 256'h17fd47fea301a90130fc92fcfcfe00f818f1a0f1e0f51bf983f5faf1a2ec20e4;
// music[4801] = 256'h97e47be1eddf1fe72bde83d60fdf9ae628e7c4d917d154cf9dc594c8dbcd3bcd;
// music[4802] = 256'h81df79f179e8fbdb34e8eff682f76ef719f599f7fcfed40054fff1f6cdf375f6;
// music[4803] = 256'hb3f2b4effcef28f686f62cefd2f18fef52ea6cf65bfe0ef74af56ff5ccf16ef4;
// music[4804] = 256'hcff0bbeeddf323f102f884f9e4ebb2f094fb6dff16fa96edf3ea59ea35ed2cf5;
// music[4805] = 256'ha5f7e1f805fbd4ff1efdf0f97e001cf606e332ddc8dc79decbde36e427e8c5dc;
// music[4806] = 256'h1adbaee73cebdce781e66ae8a6e8cee6d3e6ffe3e9e11ce78def42eeafe1aae5;
// music[4807] = 256'h85f43df052eacbeec4ec5fe5addf38dcc8db18dc9ed997d613d5b7d243d584df;
// music[4808] = 256'h0ae09ed92adab4d3c3d262df80db09d8f7df58df4ade86dc58da0ae03ae5fcdf;
// music[4809] = 256'h87db6de65ae8a8e1bae31be0f1dec5e13fe524eb8fe704e5d1e349e763ed67e2;
// music[4810] = 256'h56e1cee968e50fe362e367e335e40ee6a2ea52ee00f1d4eb67e624e5ece2e9ea;
// music[4811] = 256'h4cf551f942f85ced4be887ecfbeba3ebccef4af15ff25cf6bef389f2bef93af3;
// music[4812] = 256'h62e6cbe8bdef71f121eff7ef6af0f2eb32f0b9f466f9aaffadf072e7ffef98ef;
// music[4813] = 256'h76f223f6f2f4b4f2e4ec92f2a2f402ed90ee6bedfeeec7f2feeaa0ea8ff2cdf5;
// music[4814] = 256'h10f9e7f632edc8eccbf12eeb70e9d7f197f04deefbece8e649ed43f49aee04ee;
// music[4815] = 256'h75eebbf34d02c6026e03590c5e0b530e130df0034106e9000cfb4205f908e907;
// music[4816] = 256'hb1058802ae08c206effda7041c0d8807ee039307d505a70597072f0647097907;
// music[4817] = 256'h1008730d800185fb590536079205f5021501590206017703f30a850d6f09ac05;
// music[4818] = 256'h00059109ac0e7209f8fedeee85df07e20fe9e8e9cae98aec3cf175f08bef62ef;
// music[4819] = 256'h2aef27eec0dfbcdb98edadefc3e754e9f4e2bbdd3ae32de374e105e218e2c9e3;
// music[4820] = 256'hfbe43eeb87f503fc66f18ddda6e39af3adf92e05c70b940c860c680ad20cda0d;
// music[4821] = 256'h490b7c0893080b06c0fafaf3dcf4fff901f82defbbf460fda700c2ff29f7edf8;
// music[4822] = 256'hbffde4f99ffa030062056e0683071a0de70b1809be0d780bab035d09ed111211;
// music[4823] = 256'h7815921b1318e116081cc21d9a20f9256322cb20ac2f454015440b40f13cff3b;
// music[4824] = 256'h21410c4982484a476a49ec492a4d214e724c304e4c4e474d1c4d1f49fe470850;
// music[4825] = 256'hf952f74d514ee3508050d44baa46e5494e4cb9495549124da0503b4d314e2151;
// music[4826] = 256'h504c7d4db74cd045b840c03c0e42014456421a47fb41d74066470243d4429748;
// music[4827] = 256'hd144983ed43e503d833b503e0e397635b23aea3a993c0d3c6b36be34af30de34;
// music[4828] = 256'h6e4647506f4fc64ab847d44a054c244b414e844e494c5c489e42c545f1484d44;
// music[4829] = 256'hb4419a38432cb52d702e0c25c825322e952b4c281a2bcb27ce20fc1fa2255826;
// music[4830] = 256'h5b21a422af22d11e661e381c2e1c88208422872395217a1d2b1e881e741ae91a;
// music[4831] = 256'h7b1ae3147214d90a60fa61f806fb0a045d0a66006bfb79f77af5a4f836f1e6f1;
// music[4832] = 256'haff8b7f43bf27cf1b4f0d1ef53ef8bf13cf400f454f13ef6bdf617ec84e812e5;
// music[4833] = 256'hc9e154e6a3e9fee60ae353e250db25d5d9d815d9ebd834d3e1cacecf51d344d2;
// music[4834] = 256'h57d1afca92c9fccef6c928bfd4bb39be12c792c806bc52ba65bec0b944b666b8;
// music[4835] = 256'h93bb08bc0ac0e0c166bd24bb87b30bb2e1baa7b76bb2d9b829bf00be29ba9bb9;
// music[4836] = 256'h01ba58b731b642ba12ba98ba3ac01bbdf4b8e1bb44bdc9b915b5e6b7c1bb11bc;
// music[4837] = 256'h30bc45bf5bc914cb6ec7fbcb19cb9cc7f5c91cce31d2e9d0f2cb21cdfed12cd1;
// music[4838] = 256'h07d264d4eccfdcceead000d27ed07ec955c962cd5fd25fdc77ddc4d315d05cd7;
// music[4839] = 256'hfcd8cfd58ddcddddb6d8fbd7ebd63adb67e1cae104e085db59da4ade7fe040e2;
// music[4840] = 256'h34e247df34e259e242dae9d94bda2fdb23e371dfbade65e665e3a6eaa7f986fd;
// music[4841] = 256'h62fee6feb904ef04fdf862fa070139fdf5fd7f0286042a075b05fb01a502b400;
// music[4842] = 256'hcdfc4cfd8c036509d00308fe0904f80420fb2df8d4fc5ffdd601f0077f048f05;
// music[4843] = 256'h85054e003d074f095e0390065c070304df025f0153021d02ad0084049d06e608;
// music[4844] = 256'h4c0915f451e3cde964ea52e71ae649e689eecbef8dedafebd2ea79eec1e87cea;
// music[4845] = 256'h20f5cdefe9eb2bf17cf772ffb5001e009b07930ab9063d080105c1ff8707120a;
// music[4846] = 256'h9d03dc0077fec7fe0b04590a410d1d08dc026a053f05ac001b050c0d300e7d0a;
// music[4847] = 256'h2706460238ff14002801bc05bf0ad2062209460a200209032409d30b3706a301;
// music[4848] = 256'h610354ffaf01ab07ba07e307c1051808670863086b0bfd041e042f0745061809;
// music[4849] = 256'ha905de029d04fd05940b110fda0a2501a7ff4a066e0657078907d40540096e05;
// music[4850] = 256'h4c0079084c0f180c540a78080003cb02aa02d0079214d7070aef93eb15ebe0ea;
// music[4851] = 256'hf1f23ef742f4beef3cf3a3f53bf107f167ee24ec5eeae1e4e9e954ec8ee639eb;
// music[4852] = 256'h16edc2e260deb6e34ce29cdf4de468e2bce40feef9ef85f2daee71ec75f786fb;
// music[4853] = 256'hfcff76097e0b320ba7089c0bc20d93026ffc84f800f535047713930e3f08490f;
// music[4854] = 256'h2714bb106a0ebe0c1611e5118509a4116e1dec1b9e1dc81a6614721a0e217421;
// music[4855] = 256'hb4203b20b1257128f6214b241f2d0632d536c633142cd4288c2cbc358637ff39;
// music[4856] = 256'h263c3a35ca3a4041b53bc33ea1413e3e633f5b3f30413a45e6437c45fb3e232b;
// music[4857] = 256'hc527322b5c28112c252ace274d2b4927fa25a02b342f902d8d2e272fc1268c27;
// music[4858] = 256'h5629bc220c29962ced25ee2371237726bf283029a22d6a2b4622e81d591f9024;
// music[4859] = 256'he12a5a2ab2230b21b0216620a61e921ff8204f21462419233e1ed320a323a925;
// music[4860] = 256'hf428b0266a24481fd7190c1cdd18b418742226239f1f4c1fd51eb61ec4183b12;
// music[4861] = 256'h9313d614f4144a18cc1ae21d0622471e12166510750cde0ddb10e41158173019;
// music[4862] = 256'h7d151a174015780fd71039126b10b70ca10ce910e70fb110730ec30a46124313;
// music[4863] = 256'h70154318170e6d10e71523131912e30bbf0b2d0d7c09170b4d060201e70a7615;
// music[4864] = 256'h4413e40dd208c0ff8bfc3b0005012afce1f787fb46fe1afc49f94cfa32fe4cf8;
// music[4865] = 256'ha7f2b1f9bafa29f45cf63ff94cf6b9f4dded40eb09efe7eaf4ec83eb0de3f6e7;
// music[4866] = 256'h16e33cd987dccedb11da96d8abd0e4cbd4d2d8e14aeb72eca2e7bedfdde071ed;
// music[4867] = 256'h16f853f70cf1cbf0f8f5c1f77cf893fc5efdc5f7b1efdaecb8f158f70df66ef0;
// music[4868] = 256'h69efdeef6df2bbf48ff1edf45cf450ee62f1b8f22ef226ee9ced97f43dee29ee;
// music[4869] = 256'hd1f62ff087ed4ef2d4f0ecf08ff659f5c1ee25eefcef9ff472eec7db09dcbee2;
// music[4870] = 256'h24dc33d78ed891da61dbfcdb9cdb63dc21df9ede8ddc31dbdee05fe92fe8ece4;
// music[4871] = 256'h0de6a7e7c7e500e00ee17ce950ebe5e739e906eb11ee8eef55ea67ecabedbee7;
// music[4872] = 256'h61e985e960ea6bf021f24af0ade0e9d1f1d963dfcfda9bd9a7d70dd8bcdc78e0;
// music[4873] = 256'h6cdfa1d968d8fed8e9da4ae247e1eddce8de05dfbfdd23db5fdaa9dbc9dce2df;
// music[4874] = 256'h27df62e01de3e6e362e705e58ae224e2fbe174e61ce531e747e91ee444e94feb;
// music[4875] = 256'ha1e64eeb49f0f9ed92ea21eb7ee629e38be7c6e66fe820ed67ef74f2e2ed74ea;
// music[4876] = 256'hb6edd1ed87ebc4eac8ed54eea2eca0f041f4c2f41af2f9ebf1ecc5f47af60bf3;
// music[4877] = 256'h1cf191ef00efc0ecf8e92ef1f1f71df39ef222f6b7f2feeff6ece1e956ec0aed;
// music[4878] = 256'h48ec0cea04e886efa3f44bf0a6ed63eee3eed5edaaedd3f023f3c4f063f171f3;
// music[4879] = 256'h53ec72e93beb50e951ef9defceeae6f71907580936062f030203e4068c08aa02;
// music[4880] = 256'hf104c30e760f580d200aa404370440052406dd08050bcb0c970da1077e009703;
// music[4881] = 256'h120941074b047e046b035503cd070c083a071d0b2a0ad5069c0675062d08c508;
// music[4882] = 256'h1a055b02de005a005801d7fd06fd28030d081e0bc8fce7e3cde26fe960e6bbeb;
// music[4883] = 256'he3f39ef045ecc8e888e1d2e649f071ede4ec07ef48f183f119eb3aec9aeeaaea;
// music[4884] = 256'h32ea0eea7de73ae63ae7b8e606e3cee0b0e2b1e484e2c1e166e0cde025e7d8e7;
// music[4885] = 256'h5ae895ef00f54af022e5fbe924f8fbfe79035406cc09a00d920e880ad506ba07;
// music[4886] = 256'h6f01b5fc26fb11f4e9f13df493f96bf9ecf529faa8f6d3f45df853f709fdf3fe;
// music[4887] = 256'hcffeac01f0febaff7aff6102170ba60ad60ea615b8115f113d16de1bc6239822;
// music[4888] = 256'hca1ad21ddc238d21f321d122941fd1238d2c8f34ef3f8746e3442745cd454144;
// music[4889] = 256'h9d47214b5d4da1525e51984d774d054d9552b5561153ce4fc94af048304d3250;
// music[4890] = 256'hef5134503c4c954e1051ef49c946e74ded4d4847b7487a4cac44673f82443644;
// music[4891] = 256'h9246c94777430e4800469243f048bc45fe443143ab3eb13ecf3dda3fbf3d983b;
// music[4892] = 256'haa3d3d3a12388234623ba44f3954de4d8d4bfe4ba84d204c4e4ed954b9531750;
// music[4893] = 256'h0951504e4e4cf94d044d654cbe4afc497349bc469546eb446d49b84bfc433943;
// music[4894] = 256'hb937b02b7133d42d7322cb248629132ee429f621622271245b23ae205b231f27;
// music[4895] = 256'h32225a207f22f621b52316228922fc1f830c31034e043bffbaff02ff74fee000;
// music[4896] = 256'hfafcc3fd2a0096fa0ff664fb4904680477fe2efa7ef81af7aef772f869f138ec;
// music[4897] = 256'h40ed0ef006f2c5ed5eee79f34ef37cf3a3f028efb8f12aec79e676ea67ea9ae3;
// music[4898] = 256'h0ee363e276dba1dc22e3b0df10db27dcafd6d0d510da31d2fcd1e3d4f5cc71cc;
// music[4899] = 256'ha1c8ebc290c6e5c73cc9a8c6cac25ac2c8bfd7c104c1f7bf61c246bb3dbaeabd;
// music[4900] = 256'h38baa3baeabc93bf44bf46b9ccbb55c335c379bdb5bca3c3d6c5f9bc8bb76ec0;
// music[4901] = 256'ha0c198b7e0b904be55bcb1be87c154c2b0c259c5efc3d7c222c7f3c331c1dcc1;
// music[4902] = 256'h71c338c9bbc5ecc150c39ec44aca88cb60cd07d100ce21ca2cc8f0cc8ed1c7d0;
// music[4903] = 256'ha4cec8c93ecc85d268d17bcb19c7b4ca21d2acd5b6d1eacf4fd2f4cd41ce95d1;
// music[4904] = 256'h8cd5bddabdd520d85adba7d4dad633d688d558d7ecd4dcdbd7db31d697db1fde;
// music[4905] = 256'ha5dd63db51e221f57ef78bf409f8d3f4f9f7f6fb57f523f5a4fa68fce7fbecfa;
// music[4906] = 256'h10fcc2fdc4fc99faf8fd9f02a7ff3dfe2cff3dff12076a0b5507b708ed07a102;
// music[4907] = 256'ha5046405d9011c01d901fa04910667089b0bb60599008c00a800f703a501c301;
// music[4908] = 256'hc207ba06dc059d0311052d0af5f828e542e808edbdebc0ec8eefcaeeaee89be9;
// music[4909] = 256'he4ee99ea6ceaf8eeade98de908f08df062ef6fedf2ec98ed3cebe7e9ebe93cea;
// music[4910] = 256'hc6ebc8ee6eeca4e7bdf14b00a703ff05f509d20643ffa1ff1c037b03be07ec07;
// music[4911] = 256'he600ddff1405f804fd026506130251ff22087f071f04f9046903450444026f00;
// music[4912] = 256'he502af05cd0780047202c0025b019f010f0442064901ddfe920364020c05a00a;
// music[4913] = 256'hb0084a07ae0489008b06e90c7b057a03130a9e067d05240774048b08d1083c03;
// music[4914] = 256'h71058b08cd088109a806e003c005bb071c08f503effe93009502d4011d00a401;
// music[4915] = 256'hc40415034e04b707740a980d200c160a300adc0a68fc15e96eed27efc6ea8af3;
// music[4916] = 256'hb7f71af8baf6c5f273f03fee07ee17ec8de9b3e51de98af249ed6cebfaea1be2;
// music[4917] = 256'h00e17edd49dd18e15ddf81e66dee54f145f4cdf60df4a3ebfbee0cf563f630ff;
// music[4918] = 256'h100f08239527f61f871f611c7f19dd1725169a161011aa118815bf0ff00cc00c;
// music[4919] = 256'h0b0f0912ce0a1809ed1156134d128013fa0faa102b196d1dcf1cc71deb1e961f;
// music[4920] = 256'hd41f311e0622b529812ae029152ae92a262e102c2e2fd934eb2d9131613ae232;
// music[4921] = 256'h993183372c39ba383e2d06222225fa29db2773255c288329ba284f2ac829d029;
// music[4922] = 256'h142ac5288d26cf21f824f62be22a6a2844255e249d27dd251f258c2bf32eb729;
// music[4923] = 256'h9724e6241b28602c2b2cc22b5d2b08273e29942809263b2c45284d25762a3a28;
// music[4924] = 256'h86273f231e1f79214a1e1d2214264e205622fb26c926ff22dd1d9c1d0e1eb71e;
// music[4925] = 256'h9220a91f291e591ea721fb22a71ba517051e8a1e20183617451731170b1e8a21;
// music[4926] = 256'h471c0d1c281bc914d018eb1d841f6b21d91ae819ee1a3b15c519831ca619031c;
// music[4927] = 256'hdd1b8a1a4f18e512a11021122012a20f240f5c0ff2118315ba14281660157a0f;
// music[4928] = 256'hc510d81370142f14190e7e0daf10d20952072f0de40eef073b044b0f0a0eb403;
// music[4929] = 256'hb4083f07b402310282fe05fee7f891fae9ff11fadff85ef6c6f40bfaf2f825f7;
// music[4930] = 256'ha3f6e8f6d0f6d2f377efacea93ec47ecd8e9ffedeeeacfe59be218e189f18603;
// music[4931] = 256'hf3fdd7f271f11eeeb8ecb1f17ef13eed87e7e3e610e9f2e47ee41ae497e6aef3;
// music[4932] = 256'h7bf887f60cf3afeee4f29ff063e87cec8def2ceac2ebcef144ee2deaa9eb66e8;
// music[4933] = 256'h5ee90fed5ae940ec09edfce859ed54eb45e73ae72ae734ed0fec0cea9beacde7;
// music[4934] = 256'hd1ed3fe9c0db30dabbd91bd7c9d02ccfa3d244d3cbd8b7d699d2bcd974dd07db;
// music[4935] = 256'h19dacfde73e1f2de6dda5ed785de65df4adfbee492dc15dbc9e3cfe4c8e010dc;
// music[4936] = 256'h82e040df80da6ee1dfe231e1cae24de550e799e2f0e03ee31ae454e6b9e915e7;
// music[4937] = 256'h6ae121ead3ee49e860eb69e672d92fd55bd320d802debcdbddd948daefd910df;
// music[4938] = 256'h88e0c2d99fdee9e1c6dd63e3dde0c6deece479e443e7c5e24fdd17e580e4fee2;
// music[4939] = 256'h82e77fe9d7e841e263e127e785e91beb71ec06edb6eb3ceb44ecedeb36eccbea;
// music[4940] = 256'hf4e825e866e91dea7be889ed5beec7eaeaef41ef68f080f61ff231f264f5e6f0;
// music[4941] = 256'h83ee84f0caf141ee85ecfff168f408f0f3ed08ed25e7f9e684eb66ed55ef4aed;
// music[4942] = 256'ha8eeb4f309f227ee31eca3f128f113e86bea35ed4bea8fea77ed60ec39e80cee;
// music[4943] = 256'hc9ed19ebb7ef98e8f1e8f7ece2eba3f2e3eda6ec8feff9eb95fb5c07e0040004;
// music[4944] = 256'h8b024705a00333ffd5fea4ffea048d04ef009504810932079a03bd07140b300b;
// music[4945] = 256'h82072802cc07b20a37062b05e9014b01740625092b073a03580423073d0375fd;
// music[4946] = 256'h9a001b0855054d0364073501a0fec3026302b10571037803a6076a00cb010ffb;
// music[4947] = 256'h9aebd1ee70e8c5e38fec53e976e77ae9a8e88ee56fe6e7ecbbeabeec2eef6beb;
// music[4948] = 256'h65ef6fe703dd6de671ed80edebef0ef0e4f0daf392effdec07f20ff1e2ed6be9;
// music[4949] = 256'h98e1eee64fefe8e8ede426e741e45be5dee2cfdcc3e348e6c0e108e81ef1fff2;
// music[4950] = 256'hb7f3baf3a4e92deb6ff887f99bfff607e90a140e2a0ce50df406acffd7020afd;
// music[4951] = 256'h4dfb59fb15f850fb86f814f623f88df9caf75df5a7fa0fff4000abfe42fcdcfe;
// music[4952] = 256'h47fe2001de08b00bb80d5014061b2a1a00195718be18ac1ec51c421a1f1d0f1f;
// music[4953] = 256'h0a27db29cc2472268f2a502b752cdb2dcd31ba3c794591471f4ad24c594b5a46;
// music[4954] = 256'h1145f545f549d24cfc44f3439e47c3449746d447bc4af24c3848e348074a1b47;
// music[4955] = 256'h6e458d462b482c44cc467b4da746ed40e4435840713ebc41a740d54353460b43;
// music[4956] = 256'hce43b3417a3e913f6e428540d43ad53e103e8a3c124e575630525e558b560952;
// music[4957] = 256'hdd50a44fba4ad94d4750374cbe50c14fd347dc470f47f8458e4b144efe461944;
// music[4958] = 256'h93460b4432446f475449a2475c436444be42803eaf3b1b377d376239b73eaf3e;
// music[4959] = 256'h452a2321fc2599207f22d329a52923275623a4243723c51ef61d69122707ee04;
// music[4960] = 256'ha4059208b5014e02330cfc068702e3043b052902dbfe4d03e601bafe2f01ddff;
// music[4961] = 256'h5c03cf0232f95af8c100e008210587fd44fb7cf6a8f550f788f62cf9f4f68af0;
// music[4962] = 256'hfaefd2f38df887fab0f984f69cf2c4f3e9f386f02af125f071ec19ed3aecd9e7;
// music[4963] = 256'h8ce6dbe6f0e399dfacde11df44da33d7fddadfd84cd3d4d288d02fcf2ad046cf;
// music[4964] = 256'hd6cd5fcbbccae2c936c7bec503c43ac5c4c3f4bd2ebe84be8abcf5beddc0acbe;
// music[4965] = 256'h23bf41c271c065c085c39fc283c4cdc331be36c01cc1c3bc3bbcc2bccdbe2fc2;
// music[4966] = 256'ha1c210c2a6c00ac0abc0eebfd8c19dc38ac1b3c22dc659c68bc378c069c067c0;
// music[4967] = 256'h80bfcfc2c4c38cbf3dc29cc619c4b9c40dc885c831c8bac7cec8b9c768c655ca;
// music[4968] = 256'hb5caeac633c8eccce2cc14c92dca13ccd3ca91cbffccd5cd8fce04d177d365d1;
// music[4969] = 256'h73d0aed0b6d2c7d784d60dd4a4d2a2d8ebeeb5f6a6ef43f3fef347f320f5abf3;
// music[4970] = 256'h36f7dbf84df73ef781f75efa78f8bff6c5f9b3f827f97afce9fb1ff84df7d9f9;
// music[4971] = 256'hc4fa6bfc6bfcc6f9fcfae2fdfffd26fc9afe64ffaefac6fb6dfe08ff07fe74fb;
// music[4972] = 256'h39fe4dfed3fd9b01e0004101ab01e5fe4efe2c038f0450f37ee6c1e955e74be6;
// music[4973] = 256'h92e89ce91eed39ebd0e842eabde9ace7fae6afeaf9eb40ead5eddeefeceb82ea;
// music[4974] = 256'h20ebe8ec78f174ef1becc6ef3af05eee4aeea8f1a9f5c5f2f8f26ef4a8f1cff1;
// music[4975] = 256'h1bf192ef31ed56f39c05aa084a028204e003dd01f3012d024706a10786057506;
// music[4976] = 256'hac063005e503b1041009fb060504c606e702c101b505c703f904c00621077c09;
// music[4977] = 256'h1d0781048f06a207a904020572083b049702bb08740a0909dc079305c1058908;
// music[4978] = 256'ha2088208970a1e0a310945070706550b5b0d2809ee060c066107620979060006;
// music[4979] = 256'h52097c07e70687070305b5071a09a505ec054e08ec077104c503710324ffb4fe;
// music[4980] = 256'hf10036ffe9fc78fefcfcfbfaa8fff50004fe67f87def15eaf5e6b0e817ec43f0;
// music[4981] = 256'hcff3f4ef07f091efadebc7ed9feb37e950eb34ef65ef3be865e4a8e12fe1dce1;
// music[4982] = 256'heddcb3df08e746e816e6b9ef00052b106612d308c100840c2f12c1157f1ecc20;
// music[4983] = 256'h0d267f269721f71f301e1f1e6b1bbc1796150412e212c612230e390f58118a0c;
// music[4984] = 256'h7c0a940c0a0ccb0c39118d142e130a13f717011aa919ce19d71ab51d391d271e;
// music[4985] = 256'h0a2330244527622b67297b295a2c3d2e2f2d50218d1605176b18261af31c761f;
// music[4986] = 256'h8020501e71200523ae2286259c2825295d261c257f28c5291429f3270e272328;
// music[4987] = 256'h1a2c2d2e902b3f2d0a2db8273e28b52a872e372f332c942ea82cd129112bfe2a;
// music[4988] = 256'hc12dc02b8329f32caa29c5260c287628af2766240c2746299d2452264a28dc25;
// music[4989] = 256'ha52570225a2172255f257f23ef2231242d2674235f2130243425fc22cd21d320;
// music[4990] = 256'h421e4b1e9f1d071d9b22932332221923231d5e1cad216e21de219821e01e901d;
// music[4991] = 256'h271c661b471c7f1ccd1a0a1bce1cd01d9d1cef168217ea1b3f190e186d17db13;
// music[4992] = 256'h8e157f179313cf132816af10e310a313ee0e250f920f49112915510f450d7c0e;
// music[4993] = 256'h080bd3098808860700057204a2083b065402070182fd9d00590896064e032605;
// music[4994] = 256'h8b00bffbedf957f79bfbb9fca3fa38fdcbfa41f9f2f85df485f5ecf88ff791f7;
// music[4995] = 256'h97f9c4f715f6e0fdee089e0b0409d9061803dc00fa0100020b0060fcb1fab4fb;
// music[4996] = 256'h07fa67f6ecf356f41af424f35bf34aeeaee9c7e936e679e4f7e583e541ebeaf4;
// music[4997] = 256'h88f6dbf47ef320f078efcbf090efbcedb1ee17ef65ed64eedfebdfe88feb09ec;
// music[4998] = 256'hb2eb4ee981e8ecebf3e98eeb63e8b7d884d14dd04fceb7d0d1d4edd359d062d2;
// music[4999] = 256'hdfd10ed0e5d2fbd3aad6d7d64cd584d7b7d643d508d5a8d718d9fad470d8d9db;
// music[5000] = 256'h51d8c9d999dac0d818db79dd6cdd05df4de1e7df2adf9edee6dcf3df85e1bcde;
// music[5001] = 256'h7cde1ae064e245e3fce0e6df30e23de41ce402e542e771e91ee8e2e489e824ed;
// music[5002] = 256'h49ec7de937e796e9efe667dedbddf6dde5dcb1e096e130dfbbe06be4bfe2e6e1;
// music[5003] = 256'hf4e56ae42fe121e301e7ffe6b8e3b8e7bdea0be770e713e8f3e92aec2fe939e9;
// music[5004] = 256'h2de9c7e834eb01eabbea3eeafbe77ceeaff08eecebec06ec84ecfeede9ead7ec;
// music[5005] = 256'h04f24af076ed82ee9befbaf047f090ec32ec9aed62eb4cea86e934e8feeaf6ed;
// music[5006] = 256'ha5edd9eb1fea63ea3feac8e788e8a0ec78eb41ea8feee4eccee8bbe8d6e799eb;
// music[5007] = 256'hb7ed4dec46ee86ea72eae1eecbebf0ed4ff077ed30ed6cea11e92deaa6ebd4eb;
// music[5008] = 256'hb0ea8bf7f606a80570014a027004d0046c024702c403b2047f07dd07d0060809;
// music[5009] = 256'h4806dd036708ae08d50830071d02d70470056003f10557057c04a406c4075e05;
// music[5010] = 256'h7604f3053f03e3028503f8ffd8ffab01bc04ca051001f500a2035f024302b104;
// music[5011] = 256'h060841064803be0682fe58ecede644e7e3e7f7e895e80aea83e7b1e613e957e5;
// music[5012] = 256'h20e581ea60eb20e733e7baebdfeb8beaa8e8b9e905edcceb0fed40eef2ef97f0;
// music[5013] = 256'h90e627e256e6d7e9deed25effdf0b1f281f28ff2d9ee85ed24f0f0ebb2e36ce4;
// music[5014] = 256'h96eba6ee86eb1fe79ee619e6a4e357e2abe338e887e75de783ec1ceee4f475fb;
// music[5015] = 256'he1f1e4e692ecb5fadf01a807640c530d75108d0de109eb0e0310100b46076b03;
// music[5016] = 256'h96ffa6ff1efd42fb85ff65fc6ffbb9fe42f98efa65ff0cfe09fe38ffd303a306;
// music[5017] = 256'h0f069608620cad0f7e108f126d164917d319bd1db5208e224922f62361268925;
// music[5018] = 256'h7e25dc27612be32dbf2a122a9b2f482f6f321340ee46d34578450c44f742b644;
// music[5019] = 256'h0844674292444444d544a24878477e442f43ec45774940455443dd4495435147;
// music[5020] = 256'h274941460049f948d945be461c4794499c4991464d47f443784319446b410f4f;
// music[5021] = 256'h2a5bfb59f55d7a5c8d5726588558055a8e58e1593b5c9c5717596b59d1549856;
// music[5022] = 256'h9e53b24fbe4fea4d1c52465011490a4d9b4bf946fb491a48de46044834444f42;
// music[5023] = 256'h42423240403ffa3f943d2c3b673ecd3f5c3dcd3ae9387d3ab2394e386f397a2f;
// music[5024] = 256'h4c2597266f1da10f420f580fee0ca10cad0ac108b606bc05980680064107a809;
// music[5025] = 256'hd1090508360acb0b8707b50585059e02f1003b021503ab02a403e10165002602;
// music[5026] = 256'h18febdfa73fd5102b40601051202bbfebef72ff43ef4def2a8f0b9f20bf49af2;
// music[5027] = 256'h15f699f686f31cf3c6f068ef28f025f1adf095ed3fee99f0bbed3ae701e53ee8;
// music[5028] = 256'h5be76ae310e246e1e2e179e0bbdcf2dda6dc63d881d9a0d5b8d3cfd6fcce5ecb;
// music[5029] = 256'hb5cd3aca3fca27c96bc76ac764c55bc600c692c4bec30ac173c0b9bfc6bfafbf;
// music[5030] = 256'hd3be2cc145c177bfe3c015c29ac1e8c2c7c492c44fc57bc362c0c2c284c3dfbf;
// music[5031] = 256'hb8bf6ec2f8c185c124c22ac1ffc37fc32bbe0bc01dc28dbf91bd9dbda3bed7be;
// music[5032] = 256'h74c1acc399c264c254c4bac6e5c59cc469c52ac661c600c7a7c9c5c8c0c748cc;
// music[5033] = 256'h4acbe6c944cebfcdb9cefed21fce90cd0ed476ce3dcb9cd03cd481e1d0eb49eb;
// music[5034] = 256'hdfedc3ee44f0b7f2fcf118f3daf2d1f381f427f240f397f325f3e4f5daf58bf3;
// music[5035] = 256'h3cf451f452f3daf7d7faa0f9c3fbdbf96af6d9f9a5fb04fc4dfddafa5cfa6afd;
// music[5036] = 256'h66fdbffb94fafcf9bffc58ff4bff6dfeeffa7afbe1005200ecfd3ffc3ffc8100;
// music[5037] = 256'h8af7e3e703e78ce724e744eb23e9c9e814ec7de955ea0ceda9e9abe680e689ea;
// music[5038] = 256'h81ebe1e666ea4debe4e66febaceb85ea6ceeadebb4ea06ed1cee6df00cf0def0;
// music[5039] = 256'h0ef1f9eed2f1ccf35df014ee00efb9ee5dee56efd2ee5cf0d6f239f2cdf1a8f3;
// music[5040] = 256'h87f53ff3a6f5c501990999084805dd03dd03f104a20861099c08cd09e4099409;
// music[5041] = 256'h5807cc07ac0ddd0e550dc20ee00fca0f150fdc0ea70d270a100cac0fb90a5409;
// music[5042] = 256'h890e0e0ecb0d260fca0c000b3b0a7a0aa50a2809c209da0b580c380c3e0c0309;
// music[5043] = 256'h2605bc07dc0b0a0b1b092c0b480e130f460fef0d060e500f440b1309b60c7a0c;
// music[5044] = 256'h5409ae0bfc0b7b043c029904d9000ffda6fe610038fdf7fb2700c6ffacfc30fd;
// music[5045] = 256'h51fdd5fb03fb31fde0ff5901c30282fe9ff74df2cfe82be8eff1fdf1a3ef7df0;
// music[5046] = 256'h01efb6f095f0f5ef5ff090e968e4e2e95befaeebbef0c9fefcf9a6f3cffa00fc;
// music[5047] = 256'hf2f9dbfb40feca00c706ae0dc41187104405ae05881188120f18011e2720cf25;
// music[5048] = 256'h07223420f91fdb1aa91a3a15541131126a0db70b140d5d0b5609460a0b0abe09;
// music[5049] = 256'h290e560c7b0b71110e10430ec1115d168c184f18861c511d091fe4206611930a;
// music[5050] = 256'h6c12c70ede0da611b70feb1050124e133d15fb16dd1bb61d4d1c521c2b1e8422;
// music[5051] = 256'h3c241024f225442682258e2584242924f6263729b52ac02cf12cc42d552d2729;
// music[5052] = 256'hed295d2e292c9728112c3a2f0d2fae2f022e852c2e2e0a2d242b572cd72bb22a;
// music[5053] = 256'h7b2c802dbd2c9329c7273c29022662254029fd26ee26582a9c295b2716262526;
// music[5054] = 256'h8928e32caf2b372835295b29082bd629e7247425d126ae271e26f42391238d20;
// music[5055] = 256'h7d2354250d22b024fb21641eb9202d1de71ac41e0620341d4c1cad1eec1fac21;
// music[5056] = 256'he51f001c5c1e5b1e511bad1915174a195419ce16971bd81a831639176c12ea0f;
// music[5057] = 256'h7114ce11520dae0fdd0ee8092e0852074108c50bed0d9c0ee00c9e0bb70af108;
// music[5058] = 256'h180afb09f707d206d7042f03ff011802190026ff3408fa0fce0bb7047e002dfe;
// music[5059] = 256'hb5fe1bfddffa30fd7df966f9e0fd27f96c0435159f1358141c1420131413b70c;
// music[5060] = 256'h1f0ff50fb50ac70a6b080c09f80bad091d070c04490168ff9efdaafa6bf7dbf6;
// music[5061] = 256'h89f56ef4b4f361eec2e92be961e7c6e505e7a9e420e111e3cbe474e998f3d4f5;
// music[5062] = 256'h17f3bef32af079eccfee7ceeb6ed9cee36ebe0ea40f0baebe3d9cccec2d083d0;
// music[5063] = 256'habcda5cefdcf66cf9fcfc6d2fed2d4cfa1ce24ce35d017d218d03bcfaacf4fd2;
// music[5064] = 256'h7ed585d34ed3e5d685d6e7d311d4dcd7d0d933d75fd886d96cd685d95fdd29dc;
// music[5065] = 256'h1edcebdc03e016e0b0db93dda6dfd9dec7e17fe205df02dd31df2fe2e1e127e1;
// music[5066] = 256'hbade0adcf3de6ae1ade234e62ae619e506e50de318e5f1e956ec59ec44e9e1ea;
// music[5067] = 256'he7ef1ded29eefaf1dfe561dda4e21de15ae092e323e15ee27be473e329e33fe1;
// music[5068] = 256'hf1e320e74fe350e3ede4ece1ede207e66fe5afe61ce91ee946e906e9e0e7efea;
// music[5069] = 256'ha2ee43eabee81dee7beb88e80dea81eaeded3dee0eee85efe7ec80ed92ed3eec;
// music[5070] = 256'h87ed03ee97ed7ce977e800eafee5bbe453e564e5b1e8dbeb99eb02eb6ded88eb;
// music[5071] = 256'h0ce9dfecf0ee61ee1eec9beb0fee92eb79e9b9ebdceb80e968eb9aef49edb6ea;
// music[5072] = 256'h81ed30eed7eb60eb5fe909e8cdf64608ef077d044f056a036801b2018205b409;
// music[5073] = 256'h4a082c06f6076906a5035e033604bb078e06bd05a008d8036402a60461045507;
// music[5074] = 256'h02069f031f031701d903c20480028a0196ff80023706790249ff1200b2013602;
// music[5075] = 256'h14ff1dff1f03a80293022f046e03e8037b031bfa0eec4ae9a8eb26e8c0e7f4e7;
// music[5076] = 256'h5ce761e871e722e9a7e96ce85ee858e686e769e888e789e9a5e7a8e67feb33ea;
// music[5077] = 256'h3de5b5e8bcea50e64fe699e67ae614ea18e947e7f7e914ebc6eb25ee38ea5ae2;
// music[5078] = 256'h6fe443eafbe9abea60ed22f01bf187ee45ee99ef7cee33eb03e720e760eb63ee;
// music[5079] = 256'hc9ecaae9aaea99e72ce00be2c9e589e35ce5e6ea10edc2ee06f571fd6bfcdeef;
// music[5080] = 256'h5dedaef8e9fdc403870c440ca70f98159d12a90e090c400b050b7d06e602ed03;
// music[5081] = 256'hde03cbff0afd7dfebf012e01cefba9fb51fe82ff0d035403f1001f0290085e0d;
// music[5082] = 256'h600cd010f712e70ee111b1158b1aee1fda1f2d206d1fba21b324ab21fb231825;
// music[5083] = 256'hbd218626a12a36276127312bd228572bc9392141ca41e843f742ee439a46d745;
// music[5084] = 256'h6843ba43574728464544a847c6453e41d3437d46f4460a4a6f48cf4401496748;
// music[5085] = 256'hb443e24857495e467a5385600f60765e395ec15c4e5aaa59ce5bfb5a895a645b;
// music[5086] = 256'h9059d658c6563c559055bf533f552856f65393540e53535192540e568053e053;
// music[5087] = 256'h20538c4d574d764dbd4ac94b264a9749864b1a4a5b4954478b458c4462423e42;
// music[5088] = 256'ha4403a3f8e41df43a5427c3f9f3d4f3410265c20a6204c2140220224a11d530e;
// music[5089] = 256'h290bb510e90d110bda0d180cd105e204920842097105410493067d054f062007;
// music[5090] = 256'hdc04a008c80a5d0809071e044b010efe85fdb2ff11ff8cffc2ffd2ff4700f4fc;
// music[5091] = 256'h18fb9302230caf07d7ff92ff2cfb36f885f6c1f341f6eff4b7f445f77cf4acf3;
// music[5092] = 256'h09f343f212f3c7f304f6acf23ef14ef6b3f2a7ed01ef29edadea10ea69e699e3;
// music[5093] = 256'h2ae40be316e242e3a9e0a1dc11dc04dac1d942ddabd9b8d3e8d13bcf78d0bfd2;
// music[5094] = 256'hb2cfeaccb3cbd7cba4ca70c759c81ac9c8c523c237c13bc31bc289bf95c149c1;
// music[5095] = 256'hdbbf73c41ac4cec0b5c6e1c618c1aac395c3acbf64be58be67bf61bc93bca2c0;
// music[5096] = 256'h4abe92bd60be18be8bbefebbffbb65bd59bdb4be76bdf9bbd6bc67bd82bd0bc1;
// music[5097] = 256'h45c49bbf87bd84bfe1bfa4c438c839c9b6c903c7b4c6fcc7c7ca88cdedccadcc;
// music[5098] = 256'h0acba3d1a2e3a3ea21e663e529e82beb64ecd4e916e8ddea3eef2defc2eb62ed;
// music[5099] = 256'hc4eeecec6ff010f26bf01cf16ef273f5ebf2f1f04ff604f4e3f177f6cbf451f1;
// music[5100] = 256'hc4f274f69df7f2f56df6d3f61df7b0f84df8c2f9edfb3ffacef9eaf85af7a6f8;
// music[5101] = 256'h3cf89cf9d4f952f90dffdbf477e14de258e74de776e8f6e7bce855e9abe7c1e5;
// music[5102] = 256'h61e62de82ee772e844eaf4e9c5ea29eb1cea92e62be541e8abe832e8f1e991ea;
// music[5103] = 256'hc2e944ea36ead5e855ea5eea45e80ce9deea99ed23eeaeedb4ee7dec8fecbfee;
// music[5104] = 256'hc6ed66edd9ec27ed0def2df04af1a5f0ceef90f052f0b1ee72ef65f1a2efd0f0;
// music[5105] = 256'h3df22df06df996039a030c07f1084d0719084d07b408c609a0073909fa094808;
// music[5106] = 256'h6a086d07e507bc0a0b0b2a0b940a5c09c30b6c0cd60a240c910d270d1b0bdc0a;
// music[5107] = 256'h180ca70a8c0aeb0a90093a0a490a4509f3096d0ab009fa083709ed09dd09c909;
// music[5108] = 256'h470a7709f709be0c310c300b4d0c930af506f004bd04b8049205d005f2026f01;
// music[5109] = 256'hfe018e023102d30054019d01a3019c000fff12001aff96ffa9ff65fad7f9e1fa;
// music[5110] = 256'h4ffa69fb16fca1fd9c00f8ff92f727f814fc4feeb7eb24f212ef45f231f032f4;
// music[5111] = 256'h53054a0632037a03b5fe6cfd2e01f10390ff82fcfefa38f7f8f746f639f59df8;
// music[5112] = 256'hbef9cffc1000d903340a300e6a07dbfdd3067b109d11b11ab01d0d1dc620851e;
// music[5113] = 256'h501c321a07184918da15b613f8108a0dd40bb40a170c340c020bf70a3b0b510d;
// music[5114] = 256'h1c0d360d3f0d6d0155f762fb18fe33fda3ff4c030906ea052e07ce09e5086b0a;
// music[5115] = 256'h270e510f4d1183141917ff175b18c519c91bdd1d241e8d1e281fbe1e33212e23;
// music[5116] = 256'h6c234d247e239d249726a4251a27952a0e2bd52aed2aad295e2b502dd82af42b;
// music[5117] = 256'h9d2dfe2b282dc52b65294a2bb22b232b092bbc2a712a4229ae282529122ad029;
// music[5118] = 256'hc528d2274b260b28c329da28202a5f294e28dc29c4279a26f028ef286728aa27;
// music[5119] = 256'h6d2465231126a426492621282f293f294d295d2896264325522518255a24c623;
// music[5120] = 256'h6622242194215f22fe20001f051e951d851d951bcc1ab21c901c331d791d401c;
// music[5121] = 256'hee1eda1fc01d861d351c381ae71541111314fb15a6120f130f13d50f490f0c0e;
// music[5122] = 256'h900ce50d6c0d1e0ddd0d720d3b0ebb0ca70b1c0e130c0a0a9f0a7607c105b305;
// music[5123] = 256'h1b050107af072707fa06e00512041f025b06f80dd10d66077f03240bbf152d14;
// music[5124] = 256'hb210c211eb100510e50f390f490fe611e412df10d111bc10ea0d110f010ff70c;
// music[5125] = 256'h6c0a5509d308520546042d0416020700fbfdbbfc23f9cff5bdf4c9f25af136ee;
// music[5126] = 256'h65ec63ec31eaabe8e7e758e9c1e829e51be3b0e14de3d0df78e16cf05bf160f0;
// music[5127] = 256'ha1f0ccdd84d416d791d3ffd3cdd3dbd1c2d207d3b7d221d190d031d2e4d1e0cf;
// music[5128] = 256'hadcf4ed09ad012d28ad16ad09ad1f8d1fbd176d2ddd3c0d42cd3c9d190d1c7d3;
// music[5129] = 256'h77d591d393d3acd488d5dbd727d881d894da5bdaf4d9dfda00dc70ddbfdc7fdc;
// music[5130] = 256'h9ddd44dc57dd9fdf56debadd9bde05e1a0e132df14e01ae0e0de5ae0c1e04de2;
// music[5131] = 256'h69e3f4e24de6c8e7b7e68ee7a2e784e8ece87de9bfece5ebc3ea1aeb30e902ec;
// music[5132] = 256'h6ceef0ef92f30ceb0fe080e0d1e04ddfe8e02ee2d7e1c8e27de4aae407e466e2;
// music[5133] = 256'h17e272e36be438e566e4cbe435e7f7e763e757e77ce947eadce919eb94eb66ec;
// music[5134] = 256'h81ec9fec9eecc3e9d7ea4cec69e893e76de983e88ce675e76ce9d9e894e81cea;
// music[5135] = 256'h36eb46eb03ec09edbaeb66ea0cebc7ea17e8e1e724ea29eaaaea17eb97eabdeb;
// music[5136] = 256'h95eb28eba9ecd5ee3aed6deaefeb15eb1aec59edc6eaddf85609160854075307;
// music[5137] = 256'had04590506059f034703bd043405bd0353040504da036d067606650486041404;
// music[5138] = 256'h8902ed036205b604a104d2048005ea042402580136035b03cd00470185028a00;
// music[5139] = 256'hcd010403c8012603f302c602af03fb01b201d1014b025002110001028bfcebeb;
// music[5140] = 256'h13e686e77be666e8bfe8cfe631e665e5d0e587e6b1e6ace79ee80fe830e67ce6;
// music[5141] = 256'hade868e8a9e797e87fe836e8a5e80de8eee820ea4de826e8d3e881e755e8c9e8;
// music[5142] = 256'h5ee7eae64ae667e7dce8bee7dce76ae932ea60eaa0eb98ef36f008e97fe4c9e8;
// music[5143] = 256'hf4ec62eed5efe0effef093f277f289f1c0eee4eceaec9aea1fe769eab7ef9dea;
// music[5144] = 256'hcce79ce988e5d2e5d9e52ae40fe880e7ffe80eee6ef038f62afb2ff943f1fdf1;
// music[5145] = 256'h7efc4c0008066a0db70f4412f61099100e10140c450a1e06b103a003abff3cfe;
// music[5146] = 256'hc5fed5fc6dfb29fc16fc40fd4c00fefff1007705e007aa088e09750b130d980d;
// music[5147] = 256'h6d0e7c10f812461461158b14d713cc17ca1af71beb1c861c0c1e26205221e724;
// music[5148] = 256'h36277425a926842a7f2cc22d3030d23a9343c0402c42af433741204434445d43;
// music[5149] = 256'h08462f478a47bd46a9454845d546df454b468954a95ffc5e815f215d9f5a975b;
// music[5150] = 256'hd259c0583d594d59c4599e59b35ae05b025a3c5891587159ad59a958ab58f257;
// music[5151] = 256'h0356a35670567755eb543653d8534e538d519051fd4e7e4de14d2a4d844d2f4c;
// music[5152] = 256'hb34b164d7b4a50487248e44699454e441b436e418740c042623b0a2d72291429;
// music[5153] = 256'h0927d52757279426222666245a24302629255323c82358218c20af1c700fb40c;
// music[5154] = 256'h5211550f420ee80c540a5909f6078706af05970671066d053c068206b5050f06;
// music[5155] = 256'hdb08fb098a08e407a6055204c304440340020f0257028a033102180075ffb0ff;
// music[5156] = 256'h9704a5074302c8ff3afefcf8c0f711f6e0f47ef6e1f4e2f4a6f5bcf42cf537f4;
// music[5157] = 256'h5af452f640f6e6f564f501f4eef271f1cbee37eda1ed42edb8eb36eacbe735e5;
// music[5158] = 256'h7be397e162df08deb6dec0ded3dbd6d9aed89cd630d543d3b3d1e8d045cfd3cd;
// music[5159] = 256'h80cc97cbdeca67c9e2c71bc81dca0fca2fc8afc69bc5bcc502c506c4dac3a9c2;
// music[5160] = 256'h28c203c2cbc05ac0f9bf8bbdfebbb5bc89bc67bc7abc56bc67bde6bc07bcf4bc;
// music[5161] = 256'hdebd76becdbed6bf5fc156c202c39fc259c115c181c200c335c3e3c3fdc299c2;
// music[5162] = 256'hcfc2dbc35cc57ac553c7b7c689c9c0d8aae03fdd73de16e0e6df4ae13de12ee1;
// music[5163] = 256'h39e247e33fe428e437e434e5e8e51be669e67fe6c2e568e634e850e875e860e9;
// music[5164] = 256'h20eaa8eabdea4eebfeeb87ec4cede2edacee4fef57f076f166f14bf1f8f15cf2;
// music[5165] = 256'h7ef25bf37bf374f3e7f380f351f5b3f572f58ff77aeeffe1b4e1c9e2a4e269e3;
// music[5166] = 256'haee2a0e340e42be4dde4aee40de5e6e51ae62fe651e624e71ee816e85ae8f1e8;
// music[5167] = 256'hb6e8fee8f9e885e80ae913e916e984e981e9cae931eab5eaf3eaf8ea97ebc5eb;
// music[5168] = 256'habeb45ec0eedb0edf6ed0dee5aeeb5ee20ef3feff9eedceeb3eee7ee65ef27f0;
// music[5169] = 256'he1f006f0c5ef1ef079efb0ef1aef15ef4ef042f081f055f066f031f0e6efdef0;
// music[5170] = 256'hdeefc6f716062f087a065107bb0606082f089007b10744074b07c5060c07e107;
// music[5171] = 256'h34072e0752072c071809480acc08ef086309a4081a091109cf0822095a09e009;
// music[5172] = 256'h8409fd09020cce0c790c500c340c9a0bf70a5f0aaa0935090509b808dd07ea07;
// music[5173] = 256'h14083107ed06d206d4069a0506046f0421041904ae03d20141027d024102bc02;
// music[5174] = 256'ha2029103e3037103cc038a03c502060127ff0fffa6ff47ff14ff7bff70ffabff;
// music[5175] = 256'h3bfffcffb702fb01a7011e07620fb012310b7d04f8059207e107a20735071307;
// music[5176] = 256'h60056b034e00a1fcbcfe2105d3048dffbafdbdfa71f783f7a5f610f7fcf885fa;
// music[5177] = 256'h0ffd3e005c05600c870c5301a9fe390a1f0f8713951bf91c471f2820c41d591d;
// music[5178] = 256'h151afb179416da126811410ee10cf60ba2feb1f24ff38bf35ff3f0f4def439f6;
// music[5179] = 256'h5df759f859fa45fb47fd61ffcc000e03d3047906e808ef0bb80e581034118c12;
// music[5180] = 256'h1e14b514ea1535170f18d419ea1a071cad1dc61ee31f8320ab21f4229f23ec24;
// music[5181] = 256'h1d2635274928d02899294e2ab72a322b5c2b842b1c2c632cde2c0e2d512c542c;
// music[5182] = 256'h052c6c2ba42b182bc72adb2a792a9c2ae42ae12ae52ae82a0c2b3f2be42a612a;
// music[5183] = 256'hc42a292c2f2d302c772cb92da72c982b8729f127e82891288f28922814282728;
// music[5184] = 256'h6227a5274127f3268e2814285f2707274426fa252b250d25d9241c254a26c525;
// music[5185] = 256'h9a241c23fb21fd218b21b020b31f9e1f671f441e951d7a1c1e1c521ca61b741b;
// music[5186] = 256'h7f1a831975191819a01806169c1446174916e812cc1224120211cc102a103e10;
// music[5187] = 256'h84101b11e311a7116c119a1059107412b9126110350fb90dc00b320b7f092709;
// music[5188] = 256'h4b083e04d70b001b1e1e231b691a191edf233d21691c221b4b175914c812aa10;
// music[5189] = 256'h7710f00f650fb40f5f0f3b0fb30e590e430e780d1d0d5c0c5e0b4c0a84085707;
// music[5190] = 256'h9f05d103b702d300d0fea1fc46fa86f824f66cf3b7f1aaef67edd0ec03ec0deb;
// music[5191] = 256'h4fe9dce6ebe5eee343e4e6e0b4d171c87cc896c798c5fdc522d041d76ed483d5;
// music[5192] = 256'h1bd69ed4b4d4a0d3bed36ad398d253d2bed127d21ed200d2fad1d7d137d2d4d1;
// music[5193] = 256'h0fd292d219d2bfd1a9d1ead13dd22fd221d264d22dd3cfd322d415d586d519d5;
// music[5194] = 256'he2d59ad6e6d6d8d739d8fed8afd978d9ecd998da43db0bdbfedadcdb96db27dc;
// music[5195] = 256'h02ddc2dc5fdd8ddd2bde55df67df76e002e283e21be300e432e41ae4dce46fe5;
// music[5196] = 256'hd2e5dee66ce98eec28ec37ea4eea56ebfcebfaeba3ec6ded0cee0dee80edd1ee;
// music[5197] = 256'hccee58efa3ec5ee248e01ee34fe1abe132e2ace444e6d9e42fe6d5e5d8e61ce8;
// music[5198] = 256'h70e62ce7dfe6a2e795e894e73fe8a4e7bde8e3e98be979eacde97dea4ceb6feb;
// music[5199] = 256'h86ec87ec00ed72ec58ee7bec53e9d8f83f0792057d05c4064608ed096f084508;
// music[5200] = 256'h4d08e30782089607320753089c06d604ca040204ef05320612058b05f9016e02;
// music[5201] = 256'hb2fdc6ee80f044f7faf274f24df22bef5aee0bf229f817f9ccf7fff4d4ef6bef;
// music[5202] = 256'h1eee53ebedf095f9ebfd71fbd3f278efacefddeb27ecfcef8df457f9e5f86ff9;
// music[5203] = 256'h5cf7f2efd5ee69ee71ee6ef05bee7ff2d2f6b3f297f22bf365f060ef08efeef3;
// music[5204] = 256'h67fafff5abee77ef75f2a8f22ef1a6ee0debe2e9a4f072f8a3f90ef9c9f70ff5;
// music[5205] = 256'hc6f521f2b2e808edccf5fff610fd72fac9f4cef548eebef168f94dff4117101c;
// music[5206] = 256'hc50e2f0bba067209d907e901c709110ad506a6136d21c01eec0ff10170fbec00;
// music[5207] = 256'hc209b912701e8120ee17dd0b9304d400bcf46deb56ea50f1f6fc25f625eb25f2;
// music[5208] = 256'hf6f592f288f91c03c9fdb9f177f0daf85afd45f5ebebd2ee59f50af457f1d8f9;
// music[5209] = 256'heb016ffa4ef4fdf552f219eec1f4b805190d7c040005810e920add002907b415;
// music[5210] = 256'hcf196e1a8518e71256191b22621f8221e225c91be51b5f32d93dc73ba1337129;
// music[5211] = 256'h8d31403a29379a34732fdf377145063c26331038a535502afc28473ca94caf48;
// music[5212] = 256'h7d406d3a68352833a139044b15517d53ee5ae853304a52468052396b8f684555;
// music[5213] = 256'hb34c2455085ecb548953ba5a1961ae6757613658ff4b2047e554db5de9557240;
// music[5214] = 256'h6d37703ccb438e467d2feb1d41165911722bc1348b27d8250a1f0418290905fe;
// music[5215] = 256'h1513f3216b15ed026afcb9099d12e500f5f30dff3707990285fcc4fad0fbf0f6;
// music[5216] = 256'h08e98ee137eff3f9e6f0fbe62ceb1af4bdf1f0eeaaf0e3f530ffeaf75af0b4ef;
// music[5217] = 256'h95f2d109bb10dffc33e53ad0fcd486df79df9be72cf90b0f530a80e225c65ac7;
// music[5218] = 256'hf3d575ec38035a14fd1f551339f0cdd1f6c89dd865eb0cfe500b680ae3150d1d;
// music[5219] = 256'h640cf2029c0e182616338b35b837f23045235d1aaf1e5328d52cf32393117f11;
// music[5220] = 256'h2b1574171e2ba237be37352b2a12250ae30b0d0aeb0438fddcfe7bfdd5f98b0a;
// music[5221] = 256'h2f212b32b83ec735d11b2f0d28180b2bab23f810e614151ff120f9266e34313d;
// music[5222] = 256'hdd38462f76240b1b151b4624e428601b82131923452a13259f2c2a334323aa07;
// music[5223] = 256'h47f57ef0f0ef93f3290085094b084b0152fa13f9a0ec98d522d4a5de16df76db;
// music[5224] = 256'hd4df73e959e280d9c6df0fdf06e25aec58e909e292db0eda2ee0d3de71d671cd;
// music[5225] = 256'h8ec77bcecce4c4019e148916460abdf6afec4ef10600f60ce3064dff83033604;
// music[5226] = 256'h6e03f0fe2f03c6176f0f5ffeb10960091501750133025f0bb008ccf932f043ea;
// music[5227] = 256'hd2f14afbdefd250078ff7a05020c1d0786008200ccff1af8bcfa3805130fb91a;
// music[5228] = 256'h570ee6f776fb04065d03b6fec50a330f4efd0e0602201e201815ee0395f2b7f4;
// music[5229] = 256'h5d00350f161ad9143f15cf1ea01eaa218827f1243320771b881c5e1b31119f0a;
// music[5230] = 256'hb607e90c5a14de115713d519f91ef31f8c16fe14b51f4b215120f824fb253b27;
// music[5231] = 256'hea217217ec19f91c26198a18f81fd924b9159915b12de1388e3d81377c280329;
// music[5232] = 256'h8d2b2028bf2b91377831d217ec088d05b5126820c40f2700790c2c20f121fc15;
// music[5233] = 256'hf70c7b0c0d11ca04c5f564f3aaedc5f101f5dfebdde9cce931ed86ea5ddc25da;
// music[5234] = 256'hb9dc95dd5dea79efd4dfcadbffe6e2e6e9e0b4dc8ddd8ddda4d3b3d281daddd8;
// music[5235] = 256'h74d331d4c6d6c4d469d16cca5fc8a9d5c7e3cbe4f7d904d508d670cf3fce63d0;
// music[5236] = 256'h27cb03c7ebc9afd472e0cbdc46c583bd16d0bdd33cce7bd5e8dc44e04bd853c7;
// music[5237] = 256'h18c382ca2cd457e0aae0abd86cd8f5ce79c63dd0c8d810e60eef41e65adceccd;
// music[5238] = 256'h3acd05e39cf1dff5c8f185f99811ba14c51177120606c804b102e6eeabf15d06;
// music[5239] = 256'he80cf20e4d15521def19950c5b13b21ad2125315620ca7f769f14eec38f2f603;
// music[5240] = 256'hc70c50151121cb202e0dfefbe6f98ffb1206341213102108610b201537127211;
// music[5241] = 256'h9d19d516751217175a1c8e22f82b262c2124da1f5a1a19210f2e892a29291f30;
// music[5242] = 256'ha43900389c28e22e1f344b297b334a4243432a3d00342e3432353134b33c1342;
// music[5243] = 256'h243ba0376c3c203bc7354b37d636a933843a6a3ee6304d27b02b782eaa319735;
// music[5244] = 256'h74326c34a134c9274d27db2dbd27542f3145e14a8044aa41a940793efb3d4040;
// music[5245] = 256'h013f9738ee34b3344036f0355d30103440338e23c726f1314d2e2d29f727792d;
// music[5246] = 256'h46262d0c7405e5146613e7073913911213012607e808ba067d0c2d05f406930c;
// music[5247] = 256'h550cd50e8b081e06410259fa7a01c204520036009500befb3df3baf66bfdb9f7;
// music[5248] = 256'h41f2ebf0f6eeccea6ded9ff6ffeca7de45dfb4da11dad0e00dde1ad9aed576d6;
// music[5249] = 256'h3ed1dec9a4d755db6bd218d491cc0ac91dc98bc0c9c5cbc62fc3d8c879c092bf;
// music[5250] = 256'h84caa9bf3cb666bb43c089c39dbfa1bd99bf5bbc24b856b312b78dc202d123df;
// music[5251] = 256'hf4d877ce7cd0c4d594dc2bd7dad21cdb61d8a5d178d752e280dff3d4f9d739dc;
// music[5252] = 256'h89dac7d963dbe5dfd7db0ed730de9cdd1fc582b1b9c0dccf42c9d5c898cc1fcc;
// music[5253] = 256'ha1c6c8bc0cc294ce99d0f8d282d820d61ccbc6c7bcd06ed7c8d8dad4a2cff7d1;
// music[5254] = 256'hf9d472d3c8d129d23ad07ac6edbe54c72fd6b5d7efd354d371cbc5ca10d465d4;
// music[5255] = 256'h0bd4f6d508d1f0cb3ed081d9a6e259e888dc31d58fdedad699cff4dcf3e824ec;
// music[5256] = 256'hbce392e2d0f010f65def09e81dedfef4ceed18ee09fb8ffff1fba9f6fffd6a12;
// music[5257] = 256'haf15ed0e0f15c616b1182e288c30aa2e402d582ea52ffa2f32353238a337ab35;
// music[5258] = 256'he8339940e5436538bf404546793e1d40ce3ff53d7040293f053fa5438f40352f;
// music[5259] = 256'he727da31d3347c2f312a0f2a7c2f14317c32d032012f10362f3f7f3858325335;
// music[5260] = 256'hc03cd545433ecd343b3a8f390f3fa447b93e04441f5017434437be3a103b403c;
// music[5261] = 256'hbc425b43253fac3b023deb40b43fc03f583e1c3abb3d6446e14451348830fb3c;
// music[5262] = 256'h7e430b49684bf649b73f4a322f35413312349c3c7632d2265f26223193373e30;
// music[5263] = 256'h5231752d7f28db2d5e2f2c2f7c281f24032a4030792fb2285234603b8f33ac3b;
// music[5264] = 256'hd33ba8392f42aa3c9936b4322d2f1f344839163ca230a5221429fd287c1cb624;
// music[5265] = 256'h4c34da2e97296b30962fbc22a10de0fe7a02c1060b057f0bfa14340deafe2f00;
// music[5266] = 256'h5e0348035705f501b2fc1ef53af72403d00068051c0d9d00f5fb56f9b5f380fb;
// music[5267] = 256'h67fd85fbecfc32fa88f71cf06bed16f5d7f3a1ed25f172f632f33eee48eff7ef;
// music[5268] = 256'h4cea8de4aae4c2e49ae475e731e53ee058dedadb1fde64e23de0d3ddeedb3cd7;
// music[5269] = 256'h33d24dd46adc63d87ed203d917d7b8cd47ccf7d173dbc4da59cdaac776ce06d3;
// music[5270] = 256'h72d0f3c6a5c382d70ce745e2cedfb9e323e7bde052d627d65bda6add19da88d8;
// music[5271] = 256'h5bda00da0be0fbde0fda92dbead7f6d853d881cf43ca01cee3d32ec72ebcb0c2;
// music[5272] = 256'h87c5e1c5c3bb44b068b815be92b480abc6b1eabe42c18ec15ec779caabc5d7ba;
// music[5273] = 256'hcfb39ebbfbc778c82fc543c068b9c4bdb2c5d9c4dcbe07c0c7c8adc5f7bd2dbe;
// music[5274] = 256'hf5bf74c528c278b929be6ac156c2dec73dcb82c9b3bc1eb6debc43c34cc9afc7;
// music[5275] = 256'hbdc204c00bbc3cc0bcc6d7c67ac0a8bc03bfccbf62c221bdb1b707c1ebc005b9;
// music[5276] = 256'h3ebbd6c25ac27bbfeec87fc573b628b6d9b576bd45d63edfccd827dd12e330e3;
// music[5277] = 256'h8adc78cc8ed04fe053e085e4d4e42adaabd822d9f3d8f8dbb8e0b7e604e365dd;
// music[5278] = 256'h07e32fe4f5e0f9de0cd39ac8fec5ebc950d66adca8de89df4fdc8ade40e714ec;
// music[5279] = 256'h83e7ddeb45ec17de5ce33dea8ee870ebcbea80f075f1a2ed8af44af3e1e70be8;
// music[5280] = 256'h8bf53bf617f78afffff9e2fa56f8b0ebd8f0daf6bbfb8affb5f80ef8ebfd4bfa;
// music[5281] = 256'h43f45cf9e7fd5bffbc025a01c6035a06f804ab017c03a30d070831ffb8096715;
// music[5282] = 256'h8117f112a00f950c480bcb0bc00b2610fa138f1917188211ee12c80f3613fd11;
// music[5283] = 256'h480f202be23929318a2f132cca238e22e5318739473472352e2ea92788284f26;
// music[5284] = 256'hef2607231020722aa72daf20901e4b29ef284925361e3b0d6e0930125610600a;
// music[5285] = 256'h9d0c601021122110270f1e17be19661ac81eea174c156d1f2f1f2e181c1c7e25;
// music[5286] = 256'h352a432617198714591e7229c12f012bfd2235229b281d31932a8a1ff3218128;
// music[5287] = 256'h8e2dee2d242a7a24b424162cb5240921ca2d532b6d29222d1c24c026982d192d;
// music[5288] = 256'hb332a82d77264b2c132c2329442cf32b3b261d27182faf2c3625232561255f25;
// music[5289] = 256'h22269827022972278d2cd430e6262626cc351141b841e43ded415d487c44343e;
// music[5290] = 256'h5b3ab33b2f417c458046b1441947e5450340363fa53832314933b539923d9c3c;
// music[5291] = 256'h163c0632a91a0e0f1b18151d7b18451ef62137212c21ef19761e6f1e8916641b;
// music[5292] = 256'ha6114011f4244f233c1e531f321cda1840125c11fc14b713a3166a1d0e1bff14;
// music[5293] = 256'he7154217a015441262109a141e1a451979126c0daa0fe9153815fd0e2a0f1e14;
// music[5294] = 256'h57199616c314451abc15dc1392145b103e15971288112518ee12400f060dbd0b;
// music[5295] = 256'hde0e030c2e0ac50bc70edb0b6b06b609250cbe0aac03e902740c030561028219;
// music[5296] = 256'h4c2a4429c0241d20e3172218121c4a15e013e0120410d91cb71f61140a141a0e;
// music[5297] = 256'h8904b50b270db1068e0c720d0b09ae0b0dfe16e9bbe57ee44ee6bfed3cea1be4;
// music[5298] = 256'h65e233e24ae137dd6ade5cdeb4d9bddb62deb1db9bd97be16fe6bddd56de4ae1;
// music[5299] = 256'h25d9a8d322d294d88cdb04d21cd2ead98ddacdd4fdd0dad43cd569d0b5cc64c9;
// music[5300] = 256'hb9ccf6d122ced0ccaad2a8d170cebad382d6cad3d4d792dd09d8c6ccccc925d1;
// music[5301] = 256'hacd5ecd137d1bdd677d62acea5cb8ecf1dd277d153c9cdc82cd2ccd29ecf61cc;
// music[5302] = 256'h9ccbc2c9d0c490c924c71dcb5ce4edeb92e569e418e69be8d0e488e0c7e0cfe6;
// music[5303] = 256'ha3e6a3e36ae955e49ce380e89fe2b1e493e306e159e646e6dfe22edc22dc48d6;
// music[5304] = 256'h87c603c381c179c3dec6a2c40ac683c3dcc206c1f8bd82c243c4fcc6b6c370bc;
// music[5305] = 256'h56c287c6dec6aac7c4c30dc016c168c356bff7b9edb884ba0cbb98b47fb04bb4;
// music[5306] = 256'hdcb61eb503b5eeb4aab012b434b85cb0aea74ba791b29fb719b4adb81cb242ad;
// music[5307] = 256'he0b883b720b6f5bb1bb9f0b979b7fdb247b898b5b2b460bd0abb0aba18bd09b8;
// music[5308] = 256'h8eb861be59bf4dbb46bb6ec4dec766c701c6bac181c3f6c2e7ca91de52e286de;
// music[5309] = 256'h51df3de347e848e514e055e2a5ea16e99ae605f0f0efb4effaf1daed0af344f2;
// music[5310] = 256'heeeddcf16bf55ff835f61bf7a2f02ede62dc0be240e5a4e43adeafdda8e1e1e7;
// music[5311] = 256'hd5ea7eec60f06eecbdeb73f109f1aff30d020c0204f487f7e1f663f46e0060fe;
// music[5312] = 256'h65fc4800f6fdf1ff19009a036204e401e008f205e3fc58ff4405fc07e106ce05;
// music[5313] = 256'h5c08e20af3081f083d04300591142013f707c612b71b521588102510fd10d219;
// music[5314] = 256'h6d1f8d18471578196e1ed7193814df1ce020c025dc2b41221e1cdd1e1c224c24;
// music[5315] = 256'h5a265f28c12215278d38523ee13ad741184c8046734101430a41ba486d50494e;
// music[5316] = 256'h354c964ade47034553499e4d744bb44af24b12530b54264cb54ce546893c583f;
// music[5317] = 256'hbe42dd41273ec43a934114443d3c963da844f94497439c436b4346446d4c7656;
// music[5318] = 256'hef52134cde4c7f4a684c6256d1555f50fd4d8c49914ebc565352a94b174e2353;
// music[5319] = 256'h454f794f0c53014c09537959864c5d4bae496844bf475444b94a3253b54c1e4a;
// music[5320] = 256'h874674424143254321457747b54cfd4d0e47f4428a402243c246b0463d46fc3f;
// music[5321] = 256'h423e6a400a3c843b12402e42eb3d993d1a3ed1353e43f75826540f56b7648764;
// music[5322] = 256'h465f095ed45c6d5f30644d62465d8459a256a25aea5c9d5356502f5739574154;
// music[5323] = 256'hf9515a491446d848584136379a37f23800328d2a0d29562c59306a2e6e2b6d2b;
// music[5324] = 256'hfa27f4241a265c253924b227502eeb302d26c11a9321b0284827ee26741fdf1a;
// music[5325] = 256'h3a1d4719011caa20e2192115c3135a133916aa1471118d15cb17530ddb07430f;
// music[5326] = 256'h8a0d310895080005d4061e0948051a0276f96bf92100d0fe6703870210fdad01;
// music[5327] = 256'h9eff13fda0fff9f810ecdae3dfe522e81be544e258e2e1e445e213df3fe093de;
// music[5328] = 256'hf2dc94e6c3f7eefa84f42df34bf0c9eee3eb1ce8d5ea33ec1ceb21ea05eeeced;
// music[5329] = 256'h53e7eaee13ed1adf75e17de22fe496e674dd85dc26d9fbcb9ec781c7c4c53fbe;
// music[5330] = 256'h45b67db868ba5fb763b447b4d2b8aeb8adb2f9b13fb39daf9eaecdb0bcaf72b2;
// music[5331] = 256'h63b43babfaa6c5ad85af72a708a267a481a0869f4aa84ba2d79b7f9e7e965697;
// music[5332] = 256'h4fa0b79b079a0e9eea9b70970c90ec875289868e6b900992258e088c7d8f1689;
// music[5333] = 256'h1e86268da58c2d891f8854873287878512869f898089d4868888a48896856f87;
// music[5334] = 256'h0688fc86e7864d849f84d186cb8446834390c9a191a1ac9e989da99a009ff69e;
// music[5335] = 256'h629b3998c89899a0529ca19b30a17a98f998249fa59e61a1679e519bb69b899c;
// music[5336] = 256'hafa345a21494498bca88ec86968a598deb893e8c408fba8b748c908e5d8d818f;
// music[5337] = 256'h2b920e90e38f24935f94a9958e946a913794b5977598ac9ada9b3699c998789e;
// music[5338] = 256'heb9d6e973a97b4967b98f69dc69b319e3fa4809ecd9b86a0c79fe79e74a466a9;
// music[5339] = 256'hf9a3919b0f9f6fa3599f26a175a6e3a8fcada7ab7ea758ae32afaea955aa82ae;
// music[5340] = 256'h7fb3d6b369b39bb630b6bcb4f1b666b7ecb40bb9a2bc5fb701bbdbbec6bee6d0;
// music[5341] = 256'h80dd09d93bda3bd936d909e2c0e140dd82e297e799e6cae33be189e18be3efe4;
// music[5342] = 256'hcee6d9e770e8d2ebe3f00cf14cee8cf0bceb00dc41d4b0d13dd142db05e1a3de;
// music[5343] = 256'h80e099e1c8df88e119e74fe8e3e348e7d4f1f4f69cf6bcf861fdd0fcecfdb105;
// music[5344] = 256'hb10bc80ce7087209e90c8208fd07590c9a0a8c06310b5e158f14551316175215;
// music[5345] = 256'hae199f1bb7165c1d25225e1ec91d1e1de41dbf236825801f881e7a24ff254727;
// music[5346] = 256'h562d6c300e30e8302533e83400366e375033d92eb236cc3cd03a0e3f42433141;
// music[5347] = 256'h6d3f164030444148c3460749d3593b6895684868cd66a3655169f467ee66746b;
// music[5348] = 256'h6d6df66b5e6a186cd76de06dfc7035722f6f7f705574e1728270be6e20691c60;
// music[5349] = 256'h51540a507b5366512b524c522c4b734d5c4f8c4a344cba4ff5528750f04dbe55;
// music[5350] = 256'h7d53064ee5531f53de511259b85b9c5801599e5ad3530e51ff570e58eb533f54;
// music[5351] = 256'hf455e3552f55c858e65a3d56bb54fb571457a3543155365717585e53e751a556;
// music[5352] = 256'hbc53c74fc65075508652fc5384526f52b251664fcb4c8d4c2d4f884f004fe351;
// music[5353] = 256'h5752bd4e5c5012545b50844a9d4ba0503950da4e54503e4b994e1364c76b8462;
// music[5354] = 256'he660ee64a8679c676466e1677f6923689e61855f69641f623a5f1b631363bc5c;
// music[5355] = 256'h3259525d8f5fb75bce5ad75bd153fc467b42f542ab439340953ad93bde40ec44;
// music[5356] = 256'h7e40c537b339cf36ac35a13ea53bcc386d3e5b3fbd3bb336543a1c406b3b8438;
// music[5357] = 256'h8737a02f003102384c32fd2dfd2f0f321134c02e122d96305931f331d62f1831;
// music[5358] = 256'he230082bfe29a028b3266d24f5212d222c1ead196c199f1d0b22861fed1d511f;
// music[5359] = 256'h241ff11d1b1bec17c114e811c813481afb176e1256186015380bc40f97132c11;
// music[5360] = 256'h8911da0d9d07390db11cd0223d22ba23ac203b203c22d41ea01ddf1b1918fa15;
// music[5361] = 256'hfa15f51a961860149917c411430eea110c10cd0d0306d304f10d51021eed8dec;
// music[5362] = 256'hfcf044e945e9f8ef33eab0e6c3e63ce393e131dd18db69dcaadc4addf1db00db;
// music[5363] = 256'h32d723d471d4bad297d34ad1baccaecd16d0abd26bcc4ec537ca10cbf5c577c4;
// music[5364] = 256'ha8c58fc8c1c860c589c013bd61bd8fba5eb5efb6ceba62bbbcba99b8efb79eb8;
// music[5365] = 256'h74b368afaab737c055bd90b9e4ba3fbedac010bed4bbddbc1fbd36c0a0be03b8;
// music[5366] = 256'ha5ba8bbf09bc91b592b583ba2bb9eab787b9edb50fbcd5cc06d2e5cc2accc7cf;
// music[5367] = 256'haacd84ca5accafcc08cccac872c78fcececf79ca34c9a6c83fc6fac67fca93c9;
// music[5368] = 256'h54c599c153c569ccccc195b290aed1aa3cab02af05aca2a7d0ab84af47a8eda3;
// music[5369] = 256'h6da5fca7acac3eabd5a7b4a90dac33aa5aac3fb2e1ab77a6a8a8faa576a990af;
// music[5370] = 256'hf1ae69aa95a28da09ea9adb0d8aa7daa6faee0a04f99ed9b9198e4981794708d;
// music[5371] = 256'he692229552921b961598e49010907a97cb958d8fa98fc89187936f986e9b3797;
// music[5372] = 256'hf693ae93b6932297519af0991d998b987d962996e497fa981f9b8e98bf929f91;
// music[5373] = 256'h8d925c9f5db63bc096bc53b992ba8cba10b53cb248b5cbb724bb22c156bf61b9;
// music[5374] = 256'h4ebb3ebe7cc062c1c2be9fbfa5be15c09ac816cc96cb69c1fab26eb43eb93fb9;
// music[5375] = 256'hd2ba2eb88bb3bdb44bb9c3b93eb976bb80bc29bedfbfc2c07cc482c844c974c5;
// music[5376] = 256'h8bc33fc786c67dc65ccf57cf11c9e2cf6ed294cb4dcfbcd326d2b1d1f5ced4ce;
// music[5377] = 256'h0cd3bed57ad767da3fdd2ddad2d6e6d589d25cd5c4d75ad548d7cbd800e275e6;
// music[5378] = 256'h75dd40e262e00ed87edf11def5e2acea9de43debe4e93be49ce982e2bee302ea;
// music[5379] = 256'h7de8f8eed8ec09e795eb91f265f6d3f386faae071d0bf30d4510740fae0ee10d;
// music[5380] = 256'hed0e1a0ec70f7919131c85161b183b17990fef14f91eda1d461faf239c1ef419;
// music[5381] = 256'hac1d7b201717fb064c088d12630d78080b0a6b0a7d0d120d690b51098d071c0e;
// music[5382] = 256'hce1002133a17371211140c17cb10ca11e4156317e1153316f61bff1594148f21;
// music[5383] = 256'hca1e5b195020e01e0118251c6d2425235622db22b91b341ff8258c22bf25fb24;
// music[5384] = 256'hd01df521b5226e1d3f207721d51fdf21fd1fcb21762914278523e52333223426;
// music[5385] = 256'h4b28df255a29bc2a29297d2a072aad29712d89304d2e482c6532a335c030c838;
// music[5386] = 256'hd5477f4af74c634d3a488549f34c76530f55ec4e1352eb4f7b4d3759655bd758;
// music[5387] = 256'h125ad05d7b66386311619c65dc613966bb652055184e684e1b4ca548f045be47;
// music[5388] = 256'hd04957490e49ea4a8f4c304b0249f148364d8251534f73499f48d54b774c354d;
// music[5389] = 256'h914e494e364c0f4a274bf4498149ca49614991519d50ed470f503957fd52464e;
// music[5390] = 256'h684b774a9b4bb54e604c2e46394425468e4a634b024ae9462c412d403341fe40;
// music[5391] = 256'he83d4d3dbb43554312412345f8465546c543664277403d3d893d553b633d6341;
// music[5392] = 256'hd53a613a203cf731462bbc2bcb33354378470042c941cd436d429a4048419441;
// music[5393] = 256'h9a3f693dda3ab638ad376036a638ab3b163aed3bc53c54386739e439863a3339;
// music[5394] = 256'h66279f1aa31c7d1b9e1829174016061413146119fd18a4143614ad160016ab13;
// music[5395] = 256'hc818001b3817d81502115d0e0512b0119a0daf0de31033115c0e5e0d80119d12;
// music[5396] = 256'h760d360cd10ecd0fa70aed0501085707fc065a0805063807230a8507cbff94ff;
// music[5397] = 256'hfa07a9069800fb019f03de0350066803b4fb86fce8fe45fd63ff9c01e701a300;
// music[5398] = 256'hf6fd3afb5cfa62fdeafd45ffa302fd0060fedafb25faa5f7a1fac70bee14aa11;
// music[5399] = 256'ha213121516142f154f14c91117102f10b810fe0c1c0c301260124f0e330c8c0c;
// music[5400] = 256'h5d118a0f8d0d7e10e70c170ec009f8f33aeab4ef18f34af39bf10af198f2b2f1;
// music[5401] = 256'h72ed4aeb79ebd2eee9f771f70dedf9ed5af1a3e96ae5ece823ecd5ee49eedfeb;
// music[5402] = 256'h7debbae80de64ae652e683e8a7ea63e945e823e839e7f1e5b4e7b7e75ae24ce3;
// music[5403] = 256'h42e73be4cbe1fae151e041dc76dc71e0a0dc2ad921ddb0e298e58edf16ddb4df;
// music[5404] = 256'hd4dbcada20db30db29dd4cdb17dd04de96d86dd882dd07df8cdb94daeadb8cd8;
// music[5405] = 256'h55d7a5dcb5dbf2d7dbe55df4c3f1f4f0b2f1ddef9ef024f063f271f48af131ef;
// music[5406] = 256'h46ef88f091ee02eaebe71aea1fedf5efdef23df2d1f063ed68ec55edf5dc63ce;
// music[5407] = 256'h5fcf5dcf55d331d558d0a7ce50d030d45bd102d05ad584d47dd327d375d16dd0;
// music[5408] = 256'h78cdeccd95cfdcd021d2d2cef7cf9ada02e1a8dda3ded0e0cadb41d975d9f6df;
// music[5409] = 256'hc7e33bdb7cdd8fdf3bda72deeddb3edb85e112ddccde19e161dabbdad6da7fd9;
// music[5410] = 256'habda5ddae3dd4adda2d749d68ad5d9d8b8dd4cddf4dbb1d87bd867dcd9db99db;
// music[5411] = 256'hd7df93e3d8e250e058e137e5b4e521e1e6df64dc29dcbcf14e012eff1e002dfe;
// music[5412] = 256'h86fe4203a901220168ff22fb97fc45fffafea1fd9efabefd620437ffb8fd3d05;
// music[5413] = 256'hd404e5045b065f08c802b0eaf7dfbce575e5d0e94aee2debd9e939e567dbefdc;
// music[5414] = 256'h5de379dff5dc11de5cdd80dbb6d810dcb7def4dff2e26bdfe8dd5ade22daa7da;
// music[5415] = 256'h61e1f8e3f6e087e107def3d6cedab0e011e12edeefdd8cdd6bd798da02e00fde;
// music[5416] = 256'hd7de32dc61d8c8d6ddd590d891daf7dbf9db8fdb01dbf3d709d939dbdedddbdd;
// music[5417] = 256'h84d8e5db80de12dbb0dd27dddddbbedc0bd72dd7b6dd1fda10d678dbf9dd09dd;
// music[5418] = 256'h48d9b5d692e801fafff466f03cf101f4e5f510ef4befb6f5c8f5d4f51bf31ff2;
// music[5419] = 256'h6df614f568f452f537f2e4f26cf315f3bff3a6f2f7f845f4b7de07dac0d9b7d3;
// music[5420] = 256'h8dd82edb54dbfcda44d88fde42e26ede7edabed61bda0edd53d813d7f6d920d8;
// music[5421] = 256'h12d560d6a3daa7e061e2d0df85df19dfaedd31dccbdd22de35dbd3dea4dffedc;
// music[5422] = 256'h03de3ada88dbb7de22da1bdbbddb28d6ffd46ed69ed540d5b3d773d8f7d3bcd2;
// music[5423] = 256'h32d9b0d9efd446d8bbd854d3a3d5d1d614d218d4d6d65ad322d491d7efd70dd5;
// music[5424] = 256'h84d3f3d83ed8a7d59fd762d32dd336d21ad7d6ed12f63ff5c0f7adf173f0e6f4;
// music[5425] = 256'h43f88ff8d3f6e3f676f254f22af4b1f472fb41fa1ff779fb1efbd8fa62fc63fa;
// music[5426] = 256'h82fbd6ff78f5cde116e090e5f8e2f2e2f1e392e44cea0cef36ed8ae90ce9baeb;
// music[5427] = 256'hb1ee60ed26e961e8faeabcea54e810ebb9eef5ebd5eaaaf14af4a4efcff15af4;
// music[5428] = 256'h3cf0a4f24cf852f59ced74ec0af03eee07ef4bf4c2f4c5f544f97df762f3a4f3;
// music[5429] = 256'h14f25af224f9d4f6fdf470fa2bfa94fca4fc6dfa38fea0fb9ffbf2fec9fdabfe;
// music[5430] = 256'ha1fb13012f11c914c311e511c4126b1663181814af11c813761598180016c918;
// music[5431] = 256'he42c9c358831b6321e34423677368f32a3306e36f73acd3614387d38d037a73e;
// music[5432] = 256'h403c113b533f903b2a3cd63e6e3da63f2242ca38f326ca1f712284238a21bf22;
// music[5433] = 256'h73291e2a692ad12e0b2fab2dfe286c2636298d285d2ab42ce829c92aae2c3e2a;
// music[5434] = 256'h272c132f842d632d632c1d2dfe2e052ef5335e36ec316131372e592cc52bef29;
// music[5435] = 256'h1a2ebf30a02e8c2d862d812a362cb53119251a195820cf22d121d924d5230f24;
// music[5436] = 256'hfc25d123fb1fc11efb21cc2588238f22ba258424fa247027d527302ac629a128;
// music[5437] = 256'h4b2aa72b342ac62895298125302c6d3f28423740d243da42b54327459e44eb41;
// music[5438] = 256'h1040a642be429b42e4424b43a9457b45dc4660487b478548b948ca454745664a;
// music[5439] = 256'h2b424c2fe22e1731c32a152b242d722f2c316431c432df3036308d315532c831;
// music[5440] = 256'he42e6730da31d32fe52f7a2f732fb130ad30792fbb2e512f7e2d852b892c522e;
// music[5441] = 256'he02ed12db42e5a2ee0289e2493273e2d8c2b5b2b8b2f662cff2b622c30261627;
// music[5442] = 256'h472980281d2b992bfa2ce62c4c28c629352a8e25e625362527232f268a27d526;
// music[5443] = 256'h3028b8296c29cb27292856290f29be291e2bc52aad2b902bec257c2d41409041;
// music[5444] = 256'hb63cd93d7b3fd941cd3cd23be2404e3d713d013f613e03435342e23f9e41933f;
// music[5445] = 256'h573de53db63e964088408d3e953d9a335825b5211e213923bd27ed24ea223924;
// music[5446] = 256'h37237122802381232821e720a8219920401e421dc01fb11ed91a4519cf197f1a;
// music[5447] = 256'h7017f019ae1ded19fe1828187c19cd1bda1574145d157d1314158115e2142a12;
// music[5448] = 256'hcb0f0513ea15191632127a0e270f51108e12bb11d90c960b930d790e3f0d9d0d;
// music[5449] = 256'h130fab0b1e077a08a00a37073208420c88077607d30ba80880083507c2034505;
// music[5450] = 256'hc702e10256029dfd540a6a1a381a9c177f167a14ab142015b8121d128a132c13;
// music[5451] = 256'h0e1564133a1162163e17f517f618d7126c11051383118e1145190d1faa10bf03;
// music[5452] = 256'h930565057d076f074a035d055e04ae02ba04e401dc000602fefe93fe80ff05fd;
// music[5453] = 256'h2ffb4efbc3fd93fe25fc92fa69f81ef9fbf986f582f337f221f205f5b3f31ff2;
// music[5454] = 256'hd3f072f00ef15aed8cece7eafee781ebcbea07e929ea61ea5fed84ea8ee581e7;
// music[5455] = 256'hf1e759e71ee785e5ede3f3e2d4e468e478e01ce265e62be544e38de43ce449e1;
// music[5456] = 256'h30e051e114def9dd8fe587e2a5dd88df12db71d959db77e21ff145f4e9f440f4;
// music[5457] = 256'h54eceaec0eea05e1d7de78ddf5deb6df14dd0be0f0e2b7e115e03fde39e088e0;
// music[5458] = 256'hcfdc9fded4dd3cdc91dcd7cc45c2fbc7f5c69fc71dc80ac315c419c40ec366c5;
// music[5459] = 256'h82c61dc40cc1bcc46cc7a8c416c300c1f9c049c2b7c0e3c00bc25ac242c2a3bd;
// music[5460] = 256'hf4b881bcacbf48be30c1e7c162bc91bb76bc24bbe2bc52beeabc5eba6eb9c2bb;
// music[5461] = 256'h3dbbbfba9ebc1fbbe4b96db90bbaa5ba47b777b71dba13bd3dbedcb930b904b9;
// music[5462] = 256'ha2b832bcc5bbd7bbeabac5b88ebb15bdf5bce2bb22bcfebce8b916b950ba85bc;
// music[5463] = 256'h4fba08b9bbc993d761d642d524d4cfd3cad4e2d3b5d006cf61d07ad079d6bedb;
// music[5464] = 256'h31d9cbd9efd7d2d5ded86bd7b9d5add7cfd962d8d9d5c4d2d8c538be30c2a5c0;
// music[5465] = 256'h80c105c57cc380c389c33bc6f8c88dc5e5c467c62ac6b3c751cc08d207d11dcd;
// music[5466] = 256'hb0cdffcb34c8ccc68fc776c9afc8c0c80bccf9cef6d24ad46cd479da9fdcfed8;
// music[5467] = 256'h1bdb25dea7ddfdde45dc64d6ffd7b8d98dd8e8da83db71daa5d838d60cd782d7;
// music[5468] = 256'h1cd6d5d377d536d8fdd3a3d42bd702d5a9d62dd562d2edd2a1d3a4d4d3d364d5;
// music[5469] = 256'h85d457d1e4d218d2c3d106d25cd121cfc3ce8ede45ec7eeb21eca9ec96ec7aeb;
// music[5470] = 256'h30ea72ebe1ea27ea2fea08eb68ece4ef26f20eefcef175f255ef23f271f20cf5;
// music[5471] = 256'h1ef6fcf5a0f7d4e7f4db87e091de39dc28df05e359e440e256e37ce4b6e2c7e0;
// music[5472] = 256'h6ee1e8e3fbe3eee40be757e8d6e956ea88ea93eb8aeb6ae95ee8c1e8aae8f7ea;
// music[5473] = 256'h3aed9decaced91f1bef06eed7bf514ff8cfe88009e025100fe00d6ff64ff7404;
// music[5474] = 256'h160576012d023406ac070f085b0a92099208140bf1098909240d6b0d530d6a0e;
// music[5475] = 256'hc70e4c11fd125c11041151125a10c010a7161117e016c2191417cd169d16ce15;
// music[5476] = 256'h42250134f831bb3084326831e23164328d3158314c312633dd355436a9374039;
// music[5477] = 256'h7f3819364435583a9e3cf23a0b3dc53bc73b903b772e0c2532273b28c2259d22;
// music[5478] = 256'he122122442235e25e726bb2332222c238924b72783269026a5294b1f2317441c;
// music[5479] = 256'hab1ad416ca1623165717c418531ae21a7b1a331b7a1a47194a189c171c19ec1a;
// music[5480] = 256'he5197a19c71a90194a1a041b5b181219fc19f0187b17bc17901b421b791a811b;
// music[5481] = 256'h40192119801a1d1b081c671c151dbf1c0e1c1b1b5e1b911c671da51e5c1d2e1d;
// music[5482] = 256'h481dfa1ada1bfc1c0a1fc81d781e982e0c3826363d388037ca3549349d32a233;
// music[5483] = 256'h0a3324336834ea34ac33fc33a2377836f1346e36aa351235ab35d1370e3abc3c;
// music[5484] = 256'h6233041c7916fa1ccd1d7b2215235f22f5239c215e22f720721ceb195718041a;
// music[5485] = 256'h27195716d1156c15aa166018641776122811ee13ce12e513c216b116a3160515;
// music[5486] = 256'hc515d21ad31c9319e018581a01182f19651b491ad01cd81d191e3f1f851d441f;
// music[5487] = 256'hfd21bf23f9263e278a2767285a27d6288f2a642997297a2ac92a8d2cb22b1029;
// music[5488] = 256'h7f29de280428c4292929c427b227e02506263026f522ac221221ce237b34f63c;
// music[5489] = 256'h7f39ef39b0383936ff351036d736653421323a33d832b531b331ec319a300f2e;
// music[5490] = 256'h792d962ef52e9f2f0530112fd02d64247a14090fc10f230eca0e930e5b0d880d;
// music[5491] = 256'h5c0d690e650e7e0bdc08e408a50ad409cf077e082b09dc069b030d032c04fe02;
// music[5492] = 256'h6200f1ff28018b00fffd73fc4cfc6ffa3df789f67ff71ff7a8f4d6f21ff445f4;
// music[5493] = 256'h1ef2f5f1cbf254f120f081f0c9ed82eb93ecf2ebb3eb85eb0dead4e995ea9cee;
// music[5494] = 256'h15f16def19f05bf19bf0bfee84edabeebdf0fbf0e9ee72efcbee77eca0ed7aeb;
// music[5495] = 256'hd0ed29fa82fe3bfa09fe950c8514a21184109d10f910d4118d0f780e370f3a0f;
// music[5496] = 256'ha70f40108810c91130111e101c13dc12451159142e150d14f413ec147f0dc6fc;
// music[5497] = 256'hb3f81dfc89fa5bfb95fc59fc92fa8afa4ffe88fd0ffbbcfa5bfa5cfa46fb3cfc;
// music[5498] = 256'ha7fb99fb91f9cef60bfa91fb45f9d6f9e8fb1afce3fa34fb5dfb46fa33fa11fa;
// music[5499] = 256'h91f906f87bf78ff96af954f695f438f4aff4fdf6c7f788f6a8f6c7f67df51bf3;
// music[5500] = 256'ha7f239f30af372f6dbf75bf7ecf92ff4a1e90de853eb46ed25edb3eb69ec8cee;
// music[5501] = 256'hfbecfbebc0ed66edebedb2ee00ee73ecc4eaf9ec16ecfcef0e004f05eb01c403;
// music[5502] = 256'h9703e7029a03ac03560320022b0273037e04810595061d06c8045b053507f908;
// music[5503] = 256'h21082e07cf0625060909e20002efdeeb04ee7cebb7ec76eec1ee06ef83ef8bef;
// music[5504] = 256'h3bef95ed30eaa8eca7eefeea4fec39edc0ec4cefcfed6fec39ede5ed7ef0bfef;
// music[5505] = 256'h4dedc2ec81ebffeb48ec91e92ee878e858e90dea87e7e1e51ae98deaefe879e9;
// music[5506] = 256'h30e957e7d1e79be777e724e949e700e452e303e46de555e653e739e7c0e67de9;
// music[5507] = 256'ha1ea34e903eab7eb73eb40ea02ea92ea66ecedeb7de965ea53e926e932ebe6e9;
// music[5508] = 256'h2aea87e81aee18ffd00203009d011100470189020e02e3029001780111022902;
// music[5509] = 256'h4c032b03e4025b03b7049807b208b3075c088907d9072a0b5d00e9ef7dee09ee;
// music[5510] = 256'hbfea52ebffeae4eaaaeb2cefecf0ebee32f18cef2dec27efc5ee33edc1eb5fe9;
// music[5511] = 256'h83eb8cebd7e971ebd9ec83edceecc0ec59ed9febc1eae9eaacea2fea5ce865e7;
// music[5512] = 256'h92e87fe911e916e92be927e8c2e700e8d4e9cdeb0beb20eb01ebf7e86ae7f1e4;
// music[5513] = 256'h45e680ebe9ea4ae9c2ece0edd7ec56eec4ee33ee03ef3aef51eff3ee9fee48ef;
// music[5514] = 256'h6ced67ecbced7eed54ed8dec06ee57ef5aeb27f3770472087205cf0586056004;
// music[5515] = 256'h4e046904e103360445048f04fb06b3086f08a008050bbb0b6d0bf50cb00c450d;
// music[5516] = 256'hbb0cae0b090d8a01a7f24ef253f29fef24f10cf1a5f091f8d1028403be01e802;
// music[5517] = 256'h72024c014000f4fe94fcfdfaeafcdafdfcfc17fe13004fff97fee5ffa3ff09ff;
// music[5518] = 256'h1cfebffc0dfdc2fc29fc44fb33fa01fa82f9e1f97bfac6fa99fad9f994fa79fa;
// music[5519] = 256'h82f9cef98bf9ebf7a8f62bf706f74ff6aff691f750f940fa6efa24fb12fc9efc;
// music[5520] = 256'h1efccafcbefcc4fbeafb3ffb19fbaefaa5fadbfb17fbe9f96df617f515f7aef5;
// music[5521] = 256'h74fe080ed80f270d730d420c410c6d0c390cd70c2d0c8a0b590b260b620ce60d;
// music[5522] = 256'ha21172113406cf002e0333013f02d1029002a70340f692e8e1e954ea6ce9ece9;
// music[5523] = 256'h43e981ea33ea4fe95cea52ea1cea4aea52e9f7e60de5f2e472e51de5dee471e6;
// music[5524] = 256'he1e667e5d4e473e466e5bee6bee5dce49de446e400e46fe383e285e176e1f7e1;
// music[5525] = 256'hd2e12fe120e180e192e1e4e10be229e226e16bdfa4dfcbdf64e075e116e007df;
// music[5526] = 256'hc7dfa5e1aee2ece201e434e4a2e5dde705e8c2e703e71be631e5c6e49ce4f3e3;
// music[5527] = 256'h19e4f1e3c1e31de3efe32fe4f7e186ecbffb82fcccfa7dfb6bfb5dfb4afa5ffb;
// music[5528] = 256'hdafb27fb65fbb5fa7bfafcfae0fd630180029e01eafde0fbe8fee1011e023a05;
// music[5529] = 256'h100683f8e8ebe3eb15ece9eac6ea51ea1cea25e95fe837e8f4e85ee90ce9d0e8;
// music[5530] = 256'h8ce52ee3f7e45de518e650e995ea5dea58ea20eafaec9df1cbf296f2e0f1d7ef;
// music[5531] = 256'h03ef4cee13ee86efcff0c8f2a9f4f5f5f9f76ff9befa3dfc08fe92fe03fb7df9;
// music[5532] = 256'h60fc8afdd9fde2fe3f0078015d00a2ff9d002c017201200168010a02ba012402;
// music[5533] = 256'h3a027f01e400f0ff8cff56ff29ff35fe4bfd83fd9ffb95fbfefa5bf8ec03f111;
// music[5534] = 256'h2e11e80f71103a0f940fc40e7d0e6a0ea10d670daa0c4e0d7a0ff2101b12dc12;
// music[5535] = 256'h8112ae126312bd113b138b12ef13bc13d70454faa5fcf8fb0dfbb6fb2cfc09fd;
// music[5536] = 256'h7efce0fcbafcfefb49fc23fcfcfac5f92ef90bf86cf9aefb53faf1faf2fc67fc;
// music[5537] = 256'h65fb23fb27fb6ffb2efdc4fe95fe68fd9afccefce2fbfbfb26fc8ffb5dfce5fb;
// music[5538] = 256'h35fc3cfc4efcfdfd63fa28fd6209690d780c820dd30d020e4a0f2710a00e3c0e;
// music[5539] = 256'h900f011075102511eb117812cf12d4127613fd139d133f145314fc14ae15ac14;
// music[5540] = 256'h161505146e14b21429146321da2e2c2e392d062d5d2c412dc82cbe2c252d1a2d;
// music[5541] = 256'hef2c7d2caa2d6930cd304130d832cf332b332d330133ad3426342a3547332823;
// music[5542] = 256'h4919241bdb19c8183217e816e418d5171318601832187c197018c117b917dc16;
// music[5543] = 256'h2017e916541648168b154e156015bc142a153115821575175c128e096808a309;
// music[5544] = 256'h6b08ba0716082d081d08ba088408eb08ac097708b40725080509e4086c080d09;
// music[5545] = 256'h6c09e40a2a0c4f0cf70c0c0ca40a9b0a750b130c940c410d5d0d7f0d890c1c0c;
// music[5546] = 256'hd70c500ccd0cab0cbc0ce20c440cef0c2f0bb80b680b6e0acb186e241b23a823;
// music[5547] = 256'hfb2294220e230922f022b42268229c22672373255426952649262d273929832a;
// music[5548] = 256'h972ac72a822b6a2bcc2fb02c321a2f124d14d5124a139b13c615f0174310e208;
// music[5549] = 256'h590c231158116313401562167e193918fb131f119c0ec00c280ae1074a068c04;
// music[5550] = 256'hb1036c033e031f045a06a1063e06260783065007e3086b096b0ad009b60be60f;
// music[5551] = 256'h5e10101012119311c211ba12b21311153018531af01b771e9620c32122224e24;
// music[5552] = 256'h5c27b4289b2aa82c202d942d962e8d2ea12eb52e822e1b2f7c2d892cac2c032c;
// music[5553] = 256'hea2ecf2b942a673966414b3e0f3ef63c0d3cce3be93992376e36a936f035e836;
// music[5554] = 256'h2c3829377236e5350e359b346436c2362c3543354e3337340a2fe11b4a13cf15;
// music[5555] = 256'h8715501584125310b50f090db50bf40ab109a407a105e4067108b906a704f603;
// music[5556] = 256'h4f01e7feeefe1ffe73fdaefc20fb64facdf996f8f9f684f72df81bf660f49cf2;
// music[5557] = 256'h84f13ef12defbced79ec93e9d1e7b7e757e79be622e651e5d3e4afe43de4ade3;
// music[5558] = 256'h5ce39fe3e4e2d2e110e104dfb5dfa6e246e20fe139e1e3dfc0de46df2bde40dd;
// music[5559] = 256'he1dcd6dbeddcf2dbbdda71dbb6d91adad9d7f6d840e9a4f105ee46ef38ee23ed;
// music[5560] = 256'h39f56dfcd2fb00fbbcfb12fb5cfc99fdd8fcaafc76fc89fc2cfcb7fc18fe50ff;
// music[5561] = 256'h52ff73fdf9ffb0fab3e84fe327e654e4dce4a7e41ee4a1e58de527e542e555e4;
// music[5562] = 256'hc1e2ebe3b9e44ce3afe3b7e2e1e1f4e1ccde6cdde4dd26dd93dd7cdd37dd0ede;
// music[5563] = 256'ha5dd80dd63dfd1e0cee029e0d0df31df93ded0de38dd16dc56dcbcd934d928db;
// music[5564] = 256'h46dbc2db14dc2cdc8bdce5dcc0ddb3ddcbddc6ddd3dd80de4add54dc8ddd78de;
// music[5565] = 256'h80de21df24e0f1df12e0a0e14cdff2d419cf76d281d11ed1bbd257d0b1d1f9cf;
// music[5566] = 256'h78d21ee4c4eb65e838ea47ea8ee837e9a5e8b3e8d9e9e5e8dfe933ecb9eb57ec;
// music[5567] = 256'h86ec41ecadec1aec86edd5ed38ef82f1b9efcaf1ebea06d9a7d52fd838d606d8;
// music[5568] = 256'ha2d8ccd7c9d7e9d65fd7f6d7c9d7f3d77ed778d65bd6aed640d6e4d5b4d557d5;
// music[5569] = 256'h59d414d3c9d32fd43cd3e3d32bd4ecd3afd472d5a9d7f7d84ad7b6d62fd7dfd6;
// music[5570] = 256'h25d7d3d772d725d7d9d7eed707d8ebd846d980d98cd975d9aad9c3d9cbda0ddc;
// music[5571] = 256'h42dcd7dc38dd5cdc42db3ddb4bdc90dc21ddadde1adfb3df6ce044e01ee04fe0;
// music[5572] = 256'he3e0cde066e16ae180e002e245e07ee463f5defbf3f876fac6f941f9faf911f9;
// music[5573] = 256'h91fa89fb51fbd1fd62ff26ff1a0016000f00a5001e004401b5016202c9040e06;
// music[5574] = 256'h1b0802ff67ee7fecf1eebded7fef77ef51eff6efb5eeeeeeddf040f04beefbee;
// music[5575] = 256'he5ee75ee5aeff0edd2ed0eeec8eb2fea8ae87fe8f5e921eae4eaafebdaece4ed;
// music[5576] = 256'h2aee94f090f1d1f0b9f12bf072eef7eec0eed6efa4f0a0f0f1f14bf2b8f2f3f2;
// music[5577] = 256'hd4f2b6f389f376f310f497f4edf58cf646f67af690f608f5c7f487f6bff674f7;
// music[5578] = 256'h50f88af89cf977f988f96df95df90efa4cf924fac7f986f96ffb73f89efe900f;
// music[5579] = 256'h1214fc110113d511d0118012c8110e1385131b138c15a716f215c1169a16cf16;
// music[5580] = 256'h7d18621a6b1b771ad81bcf1bd31b2e200316a0057905bb0690052e0766061407;
// music[5581] = 256'h6c0784075a0aa509030734062d05e204fe04ea026306e1102b1375107912a212;
// music[5582] = 256'hcd107b0f310f77109a10c710bf106411a013141443130a11fc0eb10f0f108710;
// music[5583] = 256'h35115610b11073117011bb12d1121912e312ba128212d712f51217146e14f913;
// music[5584] = 256'h1814ae134a1229123a13e012a813a814dd137f14731485148615c71544166c16;
// music[5585] = 256'h7b174116541587164813d61b9d2ce32c4529942ab7292d2a232a38291d2a232a;
// music[5586] = 256'hc5298a2b922c142c1e2c902b7b2b4b2b5c2b132c3e2bf02b512b502b092d4f23;
// music[5587] = 256'h1d16ab0da0053b055c077c05c105ac07d0082008d706b0057c046c042d048a03;
// music[5588] = 256'hc40287029902b201e9019d01f900bb01d400a1ff24ff48ffb00045000e002c02;
// music[5589] = 256'h8c0279002eff8bff5cff3eff4100c000f4002d0119014401c501f0016b019301;
// music[5590] = 256'he801b4019801ce00b9006101e500290113013bff61ffd000f2002e010801ff00;
// music[5591] = 256'h5b01bf002d011201b6000f02f201930224022a0170033603870b8e1a981ba219;
// music[5592] = 256'ha11a0018ba176917ae1632176716d215fd157117371892174b18f71736179b18;
// music[5593] = 256'h1118c0163d1803171e181b1af50d1c01b2fd02fc11ffec00c20159064d073006;
// music[5594] = 256'h51054f040502a2fe12fe84fce5fa05faeef705f85bf7c3f6a3f763f797f71cf8;
// music[5595] = 256'hd6f8aef781f64bf80ef889f82df956f742fb7700aefe04fd5bfd5bfccffc12fe;
// music[5596] = 256'h94fe3e008c019d020b04290508077e087f093c0b960c010da90d000fa70f1c10;
// music[5597] = 256'he00e5f0c5c0ca50cc10c8d0d5b0d0e0db80c7e0c2d0c540c2e0c7f0b820c590b;
// music[5598] = 256'hb80a320a2307f210101f051f401cd51b001b891a46199118b117e81671167316;
// music[5599] = 256'h44189a188b175617c91625155414cc135813bb14791390138c13d504bef7b7f9;
// music[5600] = 256'h11fb08faa4fa09fcabfc55fb12fbe1f925f9d7f8eef5a2f57af5fff36ef4f7f3;
// music[5601] = 256'hb8f3caf3f5f281f200f2e8f151f10ef1c6f127f047ed43ee44f161f136f187f1;
// music[5602] = 256'h00f190f104f168f09bf003f07cf015f060efa9ef3eef30effeee04efd2eec1ee;
// music[5603] = 256'h2bef54ee8cefd5eeb5ee94f8cdfe39fc69fc64fdb4fdaffe10fea4fdc5fd0dfd;
// music[5604] = 256'h1efdb5fdf8fdc2fd7afdd1fdcffd99ffabff1afe3b0a6718e917e0163f17ce15;
// music[5605] = 256'h5316c4141414f7144c14cb13341459161d18ca179c164815f81468154615b015;
// music[5606] = 256'h7f16e2141a1665145e0483f9a7fa8bfab6fc8bfed5fdb3fd0bfc67fba5fa7efa;
// music[5607] = 256'ha9fa39f89ff5faf221f261f2b0f19df1f9f05ef1c1f110f27ff232f18cf189f1;
// music[5608] = 256'hfbf01df0e2eba8ea79ec49ed11ed41ed6eee9bed6aef60ecdadfe2dc90df4bde;
// music[5609] = 256'h43df56df0edf78df78de3ade7ede27df7edf9adfb7dfb4de12dedfdc78dc1bde;
// music[5610] = 256'h8ddee2de15dfa2de61df42dfb5de4bde21dea4dfe8de65dea9dffbddd8de98dd;
// music[5611] = 256'hdddbd3e9b4f6f8f58ef5dff499f3fdf383f39cf34cf343f3cff36bf359f47af6;
// music[5612] = 256'h6af7baf6e3f5aff57ef658f6b1f5a9f69bf529f708f575e4acdbbadec4de75e2;
// music[5613] = 256'h1ae5d8e3bbe480e3ace342e520e4c1e37ce2b5e093e2ede2b5da14d481d82cdc;
// music[5614] = 256'hf8dcc0e113e43ee465e550e4b6e3dae2fbde36dc23db5ed987d7b4d646d6cbd5;
// music[5615] = 256'hedd590d568d590d619d709d81bd997d962db84dc7bdcf7dc7ce0cce6b6e8f4e7;
// music[5616] = 256'h34e97ee920eae0eae7ea64ed4bf08ef23df63cf911fb50fd39ffac01e303e504;
// music[5617] = 256'h51076d088209ea0bf20b1b0ea00dc50d901cdc278e26c1259c252127b027ad25;
// music[5618] = 256'haa25ca24b5234a239a223c239c24f025fb2510252f237a212e21152226232c22;
// music[5619] = 256'h2f24e720f00fbd07060bc90b0a0c730b820cee0d7e0bf3090d0993099d0b810a;
// music[5620] = 256'h1e07da048e0330024501e9ff04ff4effe3feacfe7efebefe51ff48ff02fed3fb;
// music[5621] = 256'hf4fdd9ffe4fc56fb26fb56fb84fa6ff9c3f9c6f71ff7bff7b8f6abf6bdf682f6;
// music[5622] = 256'h60f563f401f4ddf2c7f2c0f222f3e7f23bf26ef282f0e8ef44f170f1bdf125f2;
// music[5623] = 256'h26f3c0f230f220f268f131f26df2c4f282f470f6f0f680f5f0f639f588f62e06;
// music[5624] = 256'h3c10c30ecd0ec60e7b0d8a0d190ea60df20d690ead0e680f830f4510de0f3c16;
// music[5625] = 256'h0822f2220422232327222823fa214024df1fba0ef509c50d0b0d2c0d6d0de90d;
// music[5626] = 256'h700ff6105410aa0fb0104e10d1102b10ce0dfd0d8b0d930d440eeb0dad0ea80e;
// music[5627] = 256'ha70eb60fec0fb5107710880e5710d013911338139f129010811194125e121213;
// music[5628] = 256'hce121713af1339139513c913c713ff131714b7142e156e158615b21500170316;
// music[5629] = 256'hcd11bd10f612a413ea13f414c715a5163517b61616167e16f016b0173d18e116;
// music[5630] = 256'hf11676173a177618b517de191120fe20932003214d208520f11fdc1fa41f381f;
// music[5631] = 256'h50202620c920ee212721b7219c23dd231c23952312230d246525d4235e26c51f;
// music[5632] = 256'h4e0e990b4c0ec20b180cd70bca0bd50b5a0c2c0efb0cd60c660dfd0c5c0d600b;
// music[5633] = 256'h9209fb09d0092e09f608df08ed08ef085b08f907f6062a0571058e0795086e07;
// music[5634] = 256'ha80726089f05b1036a03d503bb034e03830403047403920397036a061707a205;
// music[5635] = 256'h63052604f903850341028102630186ffd0ff15001800160134019f01e401d200;
// music[5636] = 256'h1d014d00b3ffc3ffb1feffff97fffffe75ff34fe6fff2efdca0062113d187416;
// music[5637] = 256'hd216ee1517155414af13741375134e13a012f312ad12a01206128712f0142814;
// music[5638] = 256'hec13ad148014f713d112c5143a0d2efedffbd8fcc0fa79fb2efbedfadbfaf1f9;
// music[5639] = 256'haafa3cfcf3fbd1fae3fa57fadbf971f8e5f5e0f506f6d5f500f665f5bef5fdf5;
// music[5640] = 256'h5ff50df41ef351f35bf388f325f329f3e0f33af31ff269f069f06ef1a5f0fcf0;
// music[5641] = 256'h2ff15df0e6f09ff11ff117f055f016f013f0b1f0d2ef3bf0e7ee6bec05ee92ee;
// music[5642] = 256'hf7edb8eea9eeebeed9efa8efb4ee02efbeee53ee88ee4beea1ef42efc6ee96ef;
// music[5643] = 256'h2aeee9eec8ec90f070014d07ec048106880520054d04f7025d036e0312030f02;
// music[5644] = 256'h71022f023c019701490160029903700301039803d003aa03490591fb4aedc8eb;
// music[5645] = 256'h2cebcde99fea53ea05eb61ea70ec78ed16edcdefb8ee66eea5ee27ed3bee88ec;
// music[5646] = 256'h3eeb47ebb5ea78eb57eb32eb8bea39e959e6b4e82ef5b5fa3cf987f9def845f9;
// music[5647] = 256'h55f89df710f799f439f500f555f48cf563f503f66ef683f6d2f667f63ff612f6;
// music[5648] = 256'h76f683f629f5c0f304f3b4f3fef405f67cf6d8f684f728f806f8fff670f650f6;
// music[5649] = 256'h7af6bbf68ff787f841f75df7cbf6dbf56af790f4e7fa1f0c6010610f1311780f;
// music[5650] = 256'hed0efc0e750e1e0e480e390e520d110e7f0d600ca50c630caa0c090ca50baf0c;
// music[5651] = 256'h760d0e0d4c0d640ef604e8f6a4f475f55cf4a7f423f4b1f3eaf338f333f2fcf3;
// music[5652] = 256'ha5f096e6eee457e6bfe47fe5d0e4c1e3b6e2e0e1d4e283e281e356e3abe192e3;
// music[5653] = 256'hd4e453e415e4abe44fe532e54be616e60be546e5cae389e238e3d9e351e390e2;
// music[5654] = 256'hbce20be32fe31ae31ae306e341e346e4f5e23ee199e102e221e342e498e4b7e4;
// music[5655] = 256'ha5e47be5dce578e503e65de6dce53ee6d0e621e7cee75ee74ae7bde64fe64ae7;
// music[5656] = 256'h51e586ecf9fc010152000403c201b8006b0075ff0eff91fe24fe73fd7afd29fd;
// music[5657] = 256'h32fd78fd53fdecfd74fd10fe26008301ad01c3010c0320f9abea68e9cde9eee8;
// music[5658] = 256'h12eacde8b5e9fcead5eb1bea07e404e411e9faebb7ed6fefdfefc2efc3f013ef;
// music[5659] = 256'h43ecaaebbfeadbe9f5e7c7e687e79ae6c1e526e62ce676e680e7fee70be814e9;
// music[5660] = 256'h92e95cea41ea50e80fe85ee943ef16f51bf3fdf1d0f16aefbdef6fef66ee82ef;
// music[5661] = 256'hb8f1b5f494f61df941fc9bfd20006002d9033006e104e30346069c0630078e07;
// music[5662] = 256'h23072608a007cf0795074f07f20750053d0e8e1efa1f621e7e1f301da21d341d;
// music[5663] = 256'hd51a671aa41959189b172c17ab15361418146a13b8127b12e1110313d315b714;
// music[5664] = 256'h5014ec14fe0769faaafab9fa34fa5ffb69fa7cfaabf9e0f859f8def7caf8a5f8;
// music[5665] = 256'h10fa1dfb55fac1fafff9d1fa5dfb45f92bf8aff7aff9a0fa7df80df8baf754f8;
// music[5666] = 256'hfef8d4f8f6f9ecf9d5f9adf9a4f8c2f892f8acf858f8f5f6daf78af84bf7c8f7;
// music[5667] = 256'h67f854f77df7a0f73df811faa3f9c1f91efac8f994fb4cfb55fbf0fcd1fc46fe;
// music[5668] = 256'h1afe99fd81fe8ffcfd02a40e990ff00e76112b114211c510a910dd103e10281a;
// music[5669] = 256'h5f2700295e281a292329ca293f29b229542a572a172b3f2b6e2b932b9e2b642b;
// music[5670] = 256'h9b2b812b442ba72c3a2c492dc82f953055309324a018011a291a51191a1a9319;
// music[5671] = 256'h771936185818181825187a1926187419e91b1b1ce81bf21bbb1b6b1a1b1b401a;
// music[5672] = 256'hf718a61afe17f7164318ee160e18a61881187f19ac19d01838168815e5153516;
// music[5673] = 256'h07179f15d613561359149a14e814db1651162817bb14ee08d4021105ce05d405;
// music[5674] = 256'hb706e3069b060b07f407b30856091b0a090a1309d608b00876096f0aed0a030b;
// music[5675] = 256'h170a5e0a4009e508cf09b7086713e62011217e20cf1f331e201fa61dea1c7c1c;
// music[5676] = 256'h2f1c261d8d1cc81b711bf91b351cb71b0e1cc41c8b1dfe1ce41c261d251f291f;
// music[5677] = 256'h5d1233081d0a320aa409380a84098a096e09ea08b408310bba0c110b230a9d0a;
// music[5678] = 256'hed0bd00b250bab0a8e092a0aa80a540cbe0dbe09f5001cfb2f00f8042a06ce0b;
// music[5679] = 256'hb70d570e710f110d330ce40971074506c5030801a7fc11fba2fa31f92cfa3ef8;
// music[5680] = 256'h53f645f72af8d8fa33fca6fc3efe71fe0aff9d00d2049a0bed0c250b770c6e0b;
// music[5681] = 256'h320b930ed60f8411ae13a21510189e199b1c351e0821102355235330003d0e3d;
// music[5682] = 256'h3f3e0b3f443ebb3e143e5a3d113d803d033d7e3cfc3c563e763fe93c4c3b623a;
// music[5683] = 256'hd5378435943343356f343a34883570294d208e22e91df217a81784170b162915;
// music[5684] = 256'hba1390112b113a10cb0f620fd00d3e0fbf0e940bb309670ae00cf60a79081307;
// music[5685] = 256'h6701cbfca5fb3efbccfaabfacbfa78fa58fad5f9b7f938fa4afab5f9e0f82ff9;
// music[5686] = 256'h4cf7c2f470f458f318f323f12aeeefedaeec2fec51ec7deb7eeb47ea26e9a7e8;
// music[5687] = 256'h0ae834e7d2e530e547e46fe36ae3bfe2c8e170e1f2e049dff7de77deb0dd2ade;
// music[5688] = 256'h60dc4edc13dc03dc90e771f1e1ef1bef01ef22ed8bece9eb18ebe0ea69ea8de9;
// music[5689] = 256'he0e859e8d2e8c3ea0dedc5ec7cec21ee43ec80ec62ed79ea17ec59e727e561f5;
// music[5690] = 256'h2cfb95f6c0f80ff88bf709f897f6e8f62cf6fbf549f67cf577f55cf5d1f5b2f6;
// music[5691] = 256'h3ff65ef625f81bf8d9f66ef706f7bef5f1f343f26df368f390f292f320f4b0f4;
// music[5692] = 256'hebf45ff53cf6adf69cf76ef7eef771f8c7f59ff4fcf4f2f393f4faf5b6f5f7f5;
// music[5693] = 256'hd0f681f6a1f6e4f66af601f7fbf7d0f82ff966f88df808f908f993f955f931f9;
// music[5694] = 256'ha1f939f9a2f9e4f971f9cafa3cfbfefa7ffc0afbb0fb8106c10e9b0d2f0e8e0e;
// music[5695] = 256'hbd0c600e390dca0d7a0ecbfcaceba0ec5bed6bec33ee31ee34ee50eecdee0cef;
// music[5696] = 256'hb9efb2f010f09cf1cbecdadf93dccbdf50df18df57df6ddf8edf37df60df26df;
// music[5697] = 256'h91deaade18df1edfb5deeade43e0a4e2b9e392e2e2e144e16fe099e020e04de0;
// music[5698] = 256'h64e1ffdfaddea6df22e038e007e18be1e3e01de01ce03ee0c2e040e180e10ce1;
// music[5699] = 256'hd5de3fdf71e242e235e13de26ae256e2b5e24ce2f7e100e240e2dae288e21ce2;
// music[5700] = 256'h37e310e4f5e368e4a0e51fe6d6e561e608e678e5f8e640e762e7d2e7bce660e7;
// music[5701] = 256'hb5e581e7b0f56dfe4bfd5ffe4ffee0fd36fef0fc62fc85fbc4fbebfcb6fcf8fc;
// music[5702] = 256'h19fd99fd6ffe60feedfeb4ffb1fff6ff3300290083019cfbbaee05ec9bedd1ec;
// music[5703] = 256'hffee2eee88ee5def9eed45ef69eda5eb6ced04ec62ecb5ecdeed5cf240f31cf2;
// music[5704] = 256'he1f12df23af2e4f1b5f2b4f2bff0b7ed7beda7ee02ee05f088f11df14ff24ef2;
// music[5705] = 256'h48f2e4f252f323f4cbf3b8f34bf227ef77ef96f0f3eedeee00f080f0e7f1caf1;
// music[5706] = 256'hd7f02ef165f1daf1ddf10bf23cf258f257f3fff204f342f3e9f24cf43cf4d6f3;
// music[5707] = 256'h04f5bbf571f614f7cdf5c0f5ecf7e1f45ef8c6074b0c300b2d0c020a780bd50a;
// music[5708] = 256'h4a0a1c0c52096e0a240be309ff0b180b770b930c5f0a500b7c0c230bd10b9e0b;
// music[5709] = 256'h1d0b910d1a064bf879f6e1f742f688f7cef890f849f8dbf8daf840f9aef9cbf7;
// music[5710] = 256'hecf7e3f7bbf719fa9ffad3fa44faf6f8f2f97ff918f8fef74ff876f7c1f681f7;
// music[5711] = 256'h19f7f2f63ef817fb94fcfafae1fc4efba9fc98113620a31cc11b7f1b3e1a7a1d;
// music[5712] = 256'hf51e4f1ecd1e141fd21ed31ee01eb61e991ef81e0e20be1f2d1e3b1e4c1f8620;
// music[5713] = 256'h4220bc1eb41e1b1e391ec11fab1f6620a31f0a1e14201520ae1f8c20211fc61f;
// music[5714] = 256'he01f531e9d1e2c1e311eba1d4d1d891d8c1c1c1d4f1aa71e6731d638b9364e38;
// music[5715] = 256'hee36d6374839a238a339cc377d37d7385437b6365136bf3577362436df35e537;
// music[5716] = 256'h4e38be375c3845375d383031fa1e291a5a1e461c951981198d180b164b19d011;
// music[5717] = 256'hb6fb3ef62ef8edf5e5f7dff334f086f1e1f17ff3a2f26cf2ddf3acf243f223f3;
// music[5718] = 256'hd0f473f546f3b6f15ef0f5eee6f0c3f1c8ee01efedf05cf104f164f1b8f53df7;
// music[5719] = 256'hc8f539f667f4d8f495f4c1eebfed62f31cf9ddf8b5f145ee0df24ff42ff332f3;
// music[5720] = 256'h97f44df599f2edf1d0f5ccf627f71bf7ddf4ddf3fef11ff3ecf54ff598f4ecf4;
// music[5721] = 256'hedf4f7f08af4db0601125910790c0a0c9c11a414fd113d0fbe0be906a507bf0d;
// music[5722] = 256'hd50e890dff0fb9114712bd11670cf40a011286110d0f4214a70de000a4fce5f6;
// music[5723] = 256'ha6f38bfa6a0197fcd8f15defbef491fb1efee5fa2dfab4f945f434f5c7fdd402;
// music[5724] = 256'hc5039dfb01f02def09f1eaf30df8faf743f78aef23e810eaf0ec37f2c3f7bafa;
// music[5725] = 256'h28fb82faccfa44f53af515f7e6eee9f27ffd9dfef8019c08130e9e0a61fffafc;
// music[5726] = 256'hac03480ce11283151618f2172e16d51810170e12bf1408191519cc162c1ab91f;
// music[5727] = 256'h6e17cb0e87116c17561acb17ae1edb205314322134350b337533be30ee29d430;
// music[5728] = 256'hb337423b2141383d063329319733a936f33b183e413e1d3d253838361d359831;
// music[5729] = 256'hf235cd3bd437e12ee624741fce17430f3815cb0e2703d314361e691c46226617;
// music[5730] = 256'h9710b313350c5b082b02c7fd600399fb28f1a1f2c9f3f1f452f963fbf7ef44e2;
// music[5731] = 256'hf3e4b2e7b0e7bfee75f3f8f765fee2fe66f584eec3f82902c305610d520dac09;
// music[5732] = 256'h810cb511e412730dcf0eaa158211700d1715621c7e20001fd018961df91ff319;
// music[5733] = 256'hf51b781e9d26152fbd2f59372f33282769291a299e250426bb2af52ea831c442;
// music[5734] = 256'h1e50464853416841cf442d4c5350fc4d03485648ff50004d1343b548e14c024b;
// music[5735] = 256'ha34c534c5946a33f134bda57e454d355074e2f45bf4afb47fb3f543a87373136;
// music[5736] = 256'h2a34783ba241ca42a93f36362736b53b263bff3601363038aa344933db35f135;
// music[5737] = 256'he635ed34b2356b388d368d32c835c5398c35db353635112e4630f32ebe20d11e;
// music[5738] = 256'h83297230dd375c394433c4309f292327a82881221927d229c32357204a136c10;
// music[5739] = 256'h031c132050257227ab22a321361c86147a18351ece1dbd1d741cda1a9217e012;
// music[5740] = 256'hca135916431a3317e913aa25772f5b2c1037bf36ff299925291b3f13ab195718;
// music[5741] = 256'h32118c154f1bff199b1bcd1ef81a8d16f312041044117e0d3210b61458ff4dee;
// music[5742] = 256'h5cf399f621f9dcf530ed8cf121fe6bff54f84afca90042fc5dfda1fb33f75bf9;
// music[5743] = 256'hbaf8c8fa9f0265051703fff9e0f368fdb305bc02f9fb7bf8d9fa49f55fefebf7;
// music[5744] = 256'h51ff55037b061b0135f7d0edacecbaf64dfe9dfc1dfd0efd7ef5e6f415f412ee;
// music[5745] = 256'h7cf230f9eefb90f7ecefdef2e5f4b7f5abf7caf1f0ef44f439f646f4c1f0eff2;
// music[5746] = 256'hc8f93a01560068f47aea1ceadef49bf61ae968f4eb0d0216621c8419c8104611;
// music[5747] = 256'hef0b560ca30bf606e411a81000102219db0cfa0ba8145a0de108c108d812ea13;
// music[5748] = 256'h94030b082d070af539f4aef4c2f415f92defd8e9bbf0bff6b3f9adf2e6ed88f0;
// music[5749] = 256'h08f2f9faeffa0ce8e0e166ed27f2baf47effe6fa20ed89f202f714f571fa44fa;
// music[5750] = 256'h7bf7c2f6cff313f51af5afee9fe8f6e98ff2a9f32ef070f514f485efccf78df8;
// music[5751] = 256'h78f316f481e97ae3c1ec4cf137f4abef31e583e434e084e405f377ecd4e73aed;
// music[5752] = 256'h43e355dbfbdc99dcdfda18d831db6de2a0df01da7fdd73df71e28ef2edfc19f8;
// music[5753] = 256'hccf68efb7cf829f1f2ef5eee25f082f7e6f697f52ef375e7b5e7def22feefbe3;
// music[5754] = 256'h72e451e438e3cce3c6e6aae537d284c706c9e0bef6be04c25abd60bec4bdb7c0;
// music[5755] = 256'habc1d4c064c835c3bab5cbb254b95dbcd4b56eb601c1aec50bbe3ebb4ac370c5;
// music[5756] = 256'h0ec3cdb660b1f8c0cac4e7c5d4ca21c41ec065bac9b57ebac7bd65c091c4f8ce;
// music[5757] = 256'h8cda99da0dd42ad43adc30e029e13fe487dffbd3f8d415e0e2db1ed755e0b4e1;
// music[5758] = 256'hf6dc64dc26dd63de3fe091e343e668e8cbe404e248e413e0fdde87e0c3e1aae7;
// music[5759] = 256'hb1e733f48609ca0950045d03e000b200b106db0868ff6401c508070286009704;
// music[5760] = 256'he006360bc30b8a05fdfee604770a0309700f0e075bf2dfeef1f1c4f7e8fc88f7;
// music[5761] = 256'h40f16bedadf110fc99fb7af842fa60f4acef3ef45df40af77bfe9dfc0df821f4;
// music[5762] = 256'hebf060f038f082fba10332f5d4e746e0e0d698ddb0e4bade39e50ce937e254e5;
// music[5763] = 256'h59dee1d8a2e557e7e3e459e7d0e7e3ea07e78ee1f6e138e0cde13fe364dde6dd;
// music[5764] = 256'hffe16fdcb9db17e5d0ec01ef4be70ee04ae12ae307e7deec1cee03ea95ebdfe9;
// music[5765] = 256'ha1de8be399e926e89ef9380a31097efe7ffdc70abe049cfa150042fb58f87e03;
// music[5766] = 256'hd8085906d204e9fe1ff7def8a2fc8afebaffd9ff0105610434f685e2fed93be1;
// music[5767] = 256'h92e153dfc7e0c5ddaae329e5dcdd48e6d1f0c3f3b1f4d6ed8eea34eefbe8a3e0;
// music[5768] = 256'ha8def4e0c1eb18f4a7ed52e8f2ea9aef13f1c9e9b6e325e73dee12f1dbef78ee;
// music[5769] = 256'h1bec7befabf1c6ed63f142edd4e4a8ead4ee20f2d6f564f7a9f90cee9de351e9;
// music[5770] = 256'h91f071f1adee53f28af176e971e773e32ce6baed6dea31eaa2e88be120e70cef;
// music[5771] = 256'h8bee2bf033e83ddd89e8a5ece1e65df9b7084807ab08df087808170acd061902;
// music[5772] = 256'hff050309fd01cd0039070b0a43049cfb33fdea0168033309e40c8108dc014bf6;
// music[5773] = 256'h1ee665e3c2e6ace4c8ebb1f032ecc2ec81eaafe8c2ec1be81ee1bee46ceb81f0;
// music[5774] = 256'h93f118e97ce04ae4a6ea22ea0eef9aefb0e0e9e230ef8cec03ed2ae8e3ddcfe2;
// music[5775] = 256'h56e98eec5fedd0e7f0e5f7e820ecf2efafef44ece8ef5cee41e56bea37ee30e6;
// music[5776] = 256'h60e961f07eebc0ebaaf2bbebd7ec81f3dae423e517ed26e647ee67f0eee63fe7;
// music[5777] = 256'h18e7bfec9df293eef5eaceea61ebf0e40de457f531068c0a910a9e0b5c07f000;
// music[5778] = 256'h69ffbbfcb1fa65fd3400bc01c706320cb90b38142d244a24571c63189d193026;
// music[5779] = 256'hcc29991300006e01fd0677086c0a1d0824034e055a05a1ff12034d0baa0d3e0a;
// music[5780] = 256'hef021e009f0014ff2e0369073901ec02ba0d2109e701be01eb00c009060dc307;
// music[5781] = 256'h0e096b034c02b709cc08dd0893060e06380bca054f071d12250e0b09380d700b;
// music[5782] = 256'h610370015b04f904a106770c2a0fb007c3051a0f8f0ca5ff3bf7d5f8ff01f305;
// music[5783] = 256'h0c0c130d8800a30075064d06170cd710a30848f8e2fd4317da1c141ab6241f21;
// music[5784] = 256'h930943034905d201d809de05a2004d0d4d0835000a016102ae085401eafd2007;
// music[5785] = 256'h2f072f0bc80695ef4be280e0bde003e758e9e0e668e7b6e320e472e728e223e9;
// music[5786] = 256'hc6f1bfe710e103e251e7b2f042ee62e8c6ed96f190ead0e428ebaff07cf089f8;
// music[5787] = 256'h07f90beda2e9c5e98ce913e574e225ee41eea7ea7af350f1d9ed6bee52e91ee9;
// music[5788] = 256'hd8eaa4e85ee718e939eb60ecf2ed2df08def16ec52f102f329e5e6dba8db85de;
// music[5789] = 256'hd3e27ceae1f26bed7deafaef76ed2beb87ed85f18ceea2edfffe8d065905650a;
// music[5790] = 256'h1f085e0e9c126c0106fd17031d02540a0b0b0d018408000d2b09b411d0109c0a;
// music[5791] = 256'hc40b56032502c202bff0f8e7d2e4c9dcade4e5eb7fe846eb15f191f580ef12e2;
// music[5792] = 256'hf0e358eab0ece4f5a6f881f3a2f2e8efb3ecb6f172fa2af73ced8af3c2fc16fb;
// music[5793] = 256'hfcfc3102ba08600daf07ce04750e811612173419df1468075708df13c714fc0e;
// music[5794] = 256'hda0e011530185d11f8fe3bf395fea708570abb15dd1b6611fd08a50bfd0fb60b;
// music[5795] = 256'h11034efdeaf448f22cfa12f896f0eaedceeeecf2fae83ce69001ad11cb0b1c0a;
// music[5796] = 256'hfd08b503360a0d16fb17351c331be3132615bd10d5138e2354243a23dd264327;
// music[5797] = 256'h672c2c29d320e724031ce010051f8220db18fb1fac1d041908180617d11e4125;
// music[5798] = 256'hd724b624e4293c27cf1eec2160213725b42b2125bc2761283c248f2c402b2324;
// music[5799] = 256'h3a263029d52b8e30a5322030aa2f3f290d1dc22077293c2a742c422cd52ba22d;
// music[5800] = 256'h9d2dd62f222ed532963f6e3f1744b14d7248f33fe2352e329e3904422f47ce41;
// music[5801] = 256'hf4393037e138cc3a2c3659397a3fa43d1b3dcc379b2a632b3a47385af44fba4a;
// music[5802] = 256'hf3529f55f94af542594bbc4ff44c094faa4c3346d448ce4df34e5f4dbf435245;
// music[5803] = 256'h424ad53f76452441f7267c266d250e1a8c1e8c21b626152f0226371ff22c2831;
// music[5804] = 256'h76261121421ae919d822af207f1e8723d623dd1fa61a40171618181c901d641b;
// music[5805] = 256'h96200d22da19f91d0f22601bb61bb01ae2166118111445087605cb0aac052206;
// music[5806] = 256'h9e0bb900bc00600398fd0806fc0449ffd4074d068501eb022bfa2af36dfec301;
// music[5807] = 256'he6fa87002e0001fa53f9c1f15cedd7f17df97efd71fc9a065315fd1b9d1bb215;
// music[5808] = 256'h26173118a2107f11af15be187c1e3e1a3814d117621cda1be518301a971b2b1c;
// music[5809] = 256'hf119cd12b4116a0751fae3fda5fb94fab504c10960059bfb2af942f78df80a02;
// music[5810] = 256'ha00005fd19fbaffd4903c2f9d1f64ef84ef162f9500141fbb1f586f378f79efb;
// music[5811] = 256'h57fa22fdd0008401d9001dfb86fc7d02cafe47fc3ef859f94c018cfd30018107;
// music[5812] = 256'h0f022f052002f0f71aff6b0760013400790645fe71f7a2ffb50025028504e1fc;
// music[5813] = 256'hb6fc2bfef5fac3fd1cfeebfc91fb77f9aaf973f71e01fa0ffa0f871059132e17;
// music[5814] = 256'h061fa11f92180a1023100618db1abf1a671d7e1c4c15a218411b5713e711300f;
// music[5815] = 256'h5214ab184a065dfbc0f484f10af9c4f2e9edaaf252f64ff997f938fdbff9b9f6;
// music[5816] = 256'h6ffb08f789f973fda0f248ed31eb39e801ec74eddeecd1eaefe6fbea95e8a4dd;
// music[5817] = 256'h11e4dbecaee57fe2b6e7bdea0feb3ae7f5e3e5e5e2e425e7faed85ea22e9e7ef;
// music[5818] = 256'h14f1f8e9a0df10de23e0a3deaae0aade23d87ad7efdb71da18d598d7a6d980d6;
// music[5819] = 256'h0bd146cd3bce69c81cc790cd10c629be58cc62e2afe7cadea9d9bddd0cde6fd5;
// music[5820] = 256'hcad7a9d955d616dda3d935d628d8d2d23bd8d8d6d5d0a1d3c1cdb1d166dbc5d5;
// music[5821] = 256'h6ec849ba3eb7c4bb44beefc05ac350c1aebccdc071c3fac303c76ac0c1c515d9;
// music[5822] = 256'hd8e092e057dad9d2edd0fad5fdda72dbc1e104e07edc4be6cee135db60e258e4;
// music[5823] = 256'h5be6ebe8a3e654e25ae009e6e1e7b3e4e7e92af059ed1aeaabe8dce3dde50aec;
// music[5824] = 256'h0beea3ef75ef45f102f164eac7ec41f794f713ec88e70ce95de7e0e89eecd0f2;
// music[5825] = 256'h06f4d5f26bf717f330f297f4fbf9eb0e350e0b066c0fc90efd0dec0c94071a0d;
// music[5826] = 256'hb7159616d30ca70a330f730c3d0cba0c9a0d9f0ff50f5d138c12610958fab1f1;
// music[5827] = 256'hb4f28cf23ff3c1f15cecd7e75ce10cde50e075e1e3e05de06bdbd1dc56e4a1e1;
// music[5828] = 256'h58e120e100da1edf9ee70de45cdc17e0c7e30ddda1dfbee3c2e770ee40e8a8e3;
// music[5829] = 256'habe2f7df5fdea1df81e9c6e722e15ce4a9e4fee714e806e25ee976f46deb72e1;
// music[5830] = 256'hf6ec4eef8aeb47ee47e737e811eb74e76ee824e346e423e838e42fe494e540e7;
// music[5831] = 256'hc9e5e3e3b9e1aee043f04afd84fd68ff9501e6fc97f142f506011501c7056b09;
// music[5832] = 256'h5604ae01c9fb82f98a03ca05d7fd28fda2fa67fb660249f5b4e50ce381de98de;
// music[5833] = 256'he1df9ee0e3e1e1e048e572e7a5e50de353dd76e1fce66edf88de4ee80ee5dddf;
// music[5834] = 256'h00e574e3d6e735eecde203e13ce9bae73be37ee058e45be4dde0b9e8a0eb37e8;
// music[5835] = 256'h7bea47e89ae32ee682ebede809e40be76ee5b6e077e4e6e718ec5fed3ce776e9;
// music[5836] = 256'hffed1dec21e976e674eb07ee17ea8ceaceeb46f299f467ed7ced4feaf0e47ae7;
// music[5837] = 256'hccee69feef04d102d808fc07c104bd04f4fb75fde9077606eb09490b4d010d05;
// music[5838] = 256'he00ae80851057d000805cdff4cfafdff4eec76dfffecf8eeb5ec85e7f5dc1de0;
// music[5839] = 256'h64e939eacce6e2e4b6e6b5ee57eecfe74fec84f080ed33e563e03de5efe29ce2;
// music[5840] = 256'he8e740e3b3e41def2bec04e698e900e95aebe1f15deecceec7ebade748ef8bea;
// music[5841] = 256'hd1e6f2efcdf2c5f495f00fe7ffe4fde5edeb3df4dcf3c2f4a8fabaf4e0ebc0ee;
// music[5842] = 256'hedf315f68df1d0ea89e8efe558ea7df5c0f2fae839ed7af1a4f2f4022e131516;
// music[5843] = 256'h9911450a620730080208840a250fa5076c07e3205129ba1d331a461678127716;
// music[5844] = 256'h24221d24b11eaf1f2612d805cd06c2fe21000e08ae01e9fd9efefcfb4403c107;
// music[5845] = 256'h8fff77000d053907aa0737fdc4fc270a250f93058901b906fffc41f634fc3d01;
// music[5846] = 256'h4508c805f4041e05d002b509e709f20aa90604faec00bf07e2067e04d1ffd501;
// music[5847] = 256'h4c056d092c0b470b0107a6ffe8050107c304a40e7a13e8129f0b68026c04a705;
// music[5848] = 256'h2d010d024005ab04ba08fd09db03ad04e40a74142e1b1c1f8922a81a6119e31a;
// music[5849] = 256'he0097303ca08cc05fa09f40a17027808170d7c076a06a60154ff7dfe8e03db08;
// music[5850] = 256'h90efc1e214edafe66de60ce942e430ea9eed16e90ee6dde451e3cbe824ee8ae9;
// music[5851] = 256'he5eaaaee3bece6e878e454e856ef8eee3beb0de928e959eaa1e5f6e216eda6ee;
// music[5852] = 256'h42ea25f24ef0bbed21f0eee4b5e28feb96f01ef1a8eac4eba2ef9de9bde99cf1;
// music[5853] = 256'hf8f06fec56eda6e95ee9c1f237f3f3f3aff6bbeeeeec6eed4ee7c0e91cef3dec;
// music[5854] = 256'hdee765ea55ec3beaecf63308ad08b207e50bc40b4e095109d0069602aa06e50a;
// music[5855] = 256'h6509d0062f016cff51034408b80c660c2f08e907120c7dff6aeb9ceeaef080e7;
// music[5856] = 256'h7be9fee9a5e5b5e891eb2be9f9e42fe462e766e558e381ea47f250f4beee97e9;
// music[5857] = 256'h76e997e8f2ef13f5e9f127f31af03af019f582f516fa67fda2004f01ddfca7ff;
// music[5858] = 256'hdb064c0b2707a307a9141c192c163811b61065166c13da0ee40f5c1234148216;
// music[5859] = 256'h931c2316f5031101b509e906a606c81278149812571739162d0fb5042005a113;
// music[5860] = 256'h241c75181213d31388133510e80bbe08020a46076107b8090909dc0c8f0bd30d;
// music[5861] = 256'hc215af14d014cf18d41cf6166e061cff0b03b40ae307e0013f0a3e13be14a20f;
// music[5862] = 256'h3f0d95141c19431ac119a61c2820c11e1922ea229b2205244d20572255220820;
// music[5863] = 256'hda223a21cb2487294326bd28eb2a0f27042dfd34382f2e2d542d80241b26d029;
// music[5864] = 256'hc52a2f332c33b931df34d730962d192dbe2c002d5f2f803351324330962ffe29;
// music[5865] = 256'hc126ed2a8630d03b2648ab42073d2541c63b9b43035c6f5f8c5aed6079609359;
// music[5866] = 256'he85bb05cb2530c514655845409533d57335a4253dd4dbd520b52634cfc4d5a4a;
// music[5867] = 256'h8d3c1033f030ac31a8335533df2fe62bc02b7d3392360c2eb22b0c2d6328b623;
// music[5868] = 256'hdb23d92dd032152d5a2ad427752b252cc32418297f2ccb298727dc1fcf1cdb1f;
// music[5869] = 256'hf022e723b322c6245f2a7f2acc20971dd020de203c21901e451cd118c91a2724;
// music[5870] = 256'h6f211020241f061bbe1e1c1d29224b2bd3255e180104a3fd6b039c0200040c05;
// music[5871] = 256'hb40399030a07770edf111f16ea1aeb188d178f1b1319a4185421a11ce3157918;
// music[5872] = 256'hef16c61b0f2078187a12c917441cc6165e180415f10187faeffd74fefcfc55fc;
// music[5873] = 256'h3bfae2f6d0f942fe97fc09f653f86cffaaf9ecf504f7abf826ff3dfd6efb9500;
// music[5874] = 256'hc001b0fd4ffadffeb001a9fb0af901fdadfc8dfa32fea3fa69f723fc47ff5d02;
// music[5875] = 256'hbcfcfbf8f6fc7bf9c4fed703aafb3cfa80007c057f03d7fe0c00eb004dfe0afc;
// music[5876] = 256'h44ffa805c608da05d8fff1fc5dffef0280fe7cfaa4faebf96c09ba17f2156618;
// music[5877] = 256'hec151c16e11cdf18f01a931f691ce1198416bc18b316f90f7c15e015ae12b418;
// music[5878] = 256'h18172c14e110b0003ffaa5ffe6fdc5fd0b00c4ff98fe72fe5803c7fe5af3f0f5;
// music[5879] = 256'h04fbecf8b8f600f7e1f52ff416fde004390207febcf761f9b5fd64f880f7c1f7;
// music[5880] = 256'h04f622f715f37ef1cdf4d6f196f323fc43fbf7f8f3f851f3aef50afa70f49eee;
// music[5881] = 256'hfdeb5df1d5f878f8a2f3abee8df514fdb5f670f3b6f409ef0ce974eb1bec0be4;
// music[5882] = 256'h5ee063e314e61ee681e8e8f2a4fc8b011603a90047ffcdffa0fe8dfc6cfe0803;
// music[5883] = 256'hb600dbf803f96ffab3f279f153f6f2f643f2a4ebd3ee1ee62bd025ce6dd082cd;
// music[5884] = 256'hfecc90cd3ecfb8c8d6c127c37cc94fc8b2bc3fbf71c121be58c460c380c037bf;
// music[5885] = 256'h6bbeabc3d8c3aec4f3bf7bb77cbb08bd33bcf6bf76beb8baa7ba46bd3ebfa7be;
// music[5886] = 256'h77bd97c0dfc2c8bec7bc0fbf8ec1bbc208c191bb91bcf7c91bcef6cfdfdd76de;
// music[5887] = 256'h74dafedda6dcfbe404eedbe805e66be325e2ebe48ae3bde45be1bae505ff7504;
// music[5888] = 256'h94fd2302a4fd2dfe2f03a5fddefef401f902ed060c03abfc8403bf0818fe82fe;
// music[5889] = 256'ha6055b02ee0a8a0648ea44e3dfea83ec0eed00ec32eb0deb47ecd0ed36f337fb;
// music[5890] = 256'h4df6c8ec1ee97fe6d6e933edc7ece5ef3ff35df6dcf7b7f6f6f7c1f8eff5f9ef;
// music[5891] = 256'h84ef83f7aaf8d5f43af363ef2bf284f8cff558f5def8faf637fa46fd4af5b3f4;
// music[5892] = 256'h56fa1cfa23fd13fa6ee8aedd40e244e312e194e6bee397de49e798ea59e875ea;
// music[5893] = 256'h59e979e7e3e715e67ae1a0e8b0fc350392febc034507f5fdecfa6200bcfce9fc;
// music[5894] = 256'h06036efeeafbcffeb9fc90fd3a024a01d6fefa02dd02acf6bde7b7de2bdd2dde;
// music[5895] = 256'h7ae256e7eee508e6d8e621e67ce6b7e195e06de77be873e319e1dbe34ce6bce4;
// music[5896] = 256'h36e19cdb96d9bbe206ebd0e70ee774e861e53be871eba0ec7bec71e4a4e320e5;
// music[5897] = 256'haee07fe554e960e84eea14e9a6e8dce714e685e617e423e38de585e8fcea1eeb;
// music[5898] = 256'heeedd9eda2e887e575e010e211ea47ebaced47ed69eb8deac4e1cfecca046008;
// music[5899] = 256'h4a079704880166044004920471020c0294020701ce05bdffccfa4204eb050105;
// music[5900] = 256'hb801400077fe49ed3ee6a1e77fe4bfe89de8efe7e7e939e642e575e342e18ce4;
// music[5901] = 256'hb1e630e595e5a2ec51eda9e41ee432e65fe2bede63df9fe8c8ed2dec86f024ee;
// music[5902] = 256'h80eab5eb12e4d1e77cee81e6a3e883e9fae39fe774e79be910ef9ced64ef2ded;
// music[5903] = 256'hc9e796ec20ed8ce76be94eebd0e89fe8b6eae3eb45eccced60ed47ed0af301f1;
// music[5904] = 256'h37e8cced0bf143eb71f82c062f09c8101a08e5fe1306d9051108e808f1069f0c;
// music[5905] = 256'hc507a804d0052301c2011e01c10444060001260166f2a0e3ece915ea52e626e9;
// music[5906] = 256'h5fe8aee648ea70ec44ecd2edbde8b9e448eb51ec8de8cfe7a1e50ae60ce7c2e3;
// music[5907] = 256'h71e5cfec6ff047ed90e6aee696effbf41ef38befededc1ec66e911e84cee45f3;
// music[5908] = 256'hf4ed33ec55f03df0d6f440f739f169f5ec005208490a0c07ca0af410060dea08;
// music[5909] = 256'h2305cd042e0d760a8904e60a220c2b0a950c650b9c0ef61d892767225123a525;
// music[5910] = 256'h441d461d59245e262924801f8a1d1e1d261e3d1f7a1ea71f89200b22d421f11e;
// music[5911] = 256'h57170f0a2807ac053a005a06c30563ff8f03fd029eff37054f08130504071f08;
// music[5912] = 256'he402c80236020301f3034103820669076efe98fd930207031b01f4ff81ffecfc;
// music[5913] = 256'h56006305fa02d002680037fcd100e6041006e50505037f031a0419016efb6df4;
// music[5914] = 256'h82f030efe1ec51ecf8f0e1ee62e7c0eb9befb2ef49f482f2ecf000f440f38fed;
// music[5915] = 256'h40eea901d40f600cdc09dc08d2074708610c7f0c9a061908d50676049a078205;
// music[5916] = 256'h5e044a031607560bb60402047bffcbf297ec8de8d7edcbf1abec0fecd8e8f7e6;
// music[5917] = 256'h5eecaced5cecf9eb2dea1fecd6efbdea07e643ebbaed7ae6a7e1d6e6a1e8f5e7;
// music[5918] = 256'h4cec61eb79ea13ecf3e98eea14ed7ef19cf6c4f5feee13e8b6e70ae9f1e545e5;
// music[5919] = 256'hfbec45f571f683f688f11ce94cea2bebede966f1dbf33befdaf304f829f239ed;
// music[5920] = 256'h71ea8cec0ff2a8f433fa02f844f26201a4102c0d140ae40c970abc041206fd09;
// music[5921] = 256'h83075507b9086f051304f300aafff1071f0ae6055c044f060e08ccf89ae9d7f3;
// music[5922] = 256'h8bff89fc3ff713f5adf49df9b3fb65f523f619f853f869ff9afe92fb3f01f308;
// music[5923] = 256'h1e0f770e830e860e260c4a0fbe0f72101e118f0d8f10a110fb0d9c10aa123010;
// music[5924] = 256'habff1efad90ad70a790616105d15571adc19440f590b600d0d098f01c600d8fe;
// music[5925] = 256'hbffaa0fd3ffceef5dbf3e1f1caf0ccf2bbf3f6f503fcc5fb6ff610fc6f0c6517;
// music[5926] = 256'hd915bf17fb1f2e2151226a238320d5225527be2a732f9d2e622c72333e35292f;
// music[5927] = 256'h57308232f133c42d862215212e1f4d236426991f50240826ab28092ff1283329;
// music[5928] = 256'h9f299829482de52691291b2ecf2a612bb22a562f8b33802c6d270a2a562ddb2b;
// music[5929] = 256'hb32add293e29ae2d902f2d2f19345335bb2cd127e62d3a3516370633242e3e2e;
// music[5930] = 256'h083002305436724205450445a548ee4702482241c836cf3ade3fa93ed83e5540;
// music[5931] = 256'h52438243843ad9354048375bcf57cb53c858ea59bb56bc531c5127531e57fe53;
// music[5932] = 256'hf44e884ab5485d4c214b164c6a4f9a4a99492742ae2e8e2c7531b629fe28ba2b;
// music[5933] = 256'he225bc253727f627f82b94290c27f8243c1f8a1e4421d4249923f820df22b21d;
// music[5934] = 256'hb21b92211d2004210224431e021cc01e2e1b66180b1d441f461bf61ac920df1f;
// music[5935] = 256'ha81848155e188821e61e1d14b418031e701b8710d50095007b03750449088e05;
// music[5936] = 256'h2107b906ee02ec04ad05410b7d0858ff9e02f7fe64ff8c110e1d1e1eb41ced1c;
// music[5937] = 256'hf61eb3216a2092176e17a9203f215c184414ad1aea194814671822186d15af1c;
// music[5938] = 256'hfb168800cefa9bffb5fb18fda1fdbefa90fcdffa42ff5901f8f7bef668f73bf9;
// music[5939] = 256'h50ff92fedc0031038cfd58fafefb180056031d02edfc08f7c2f747fe2efe4af7;
// music[5940] = 256'hcaf712fed502220346005b028bffcefc54044d02ed0020039efd8a02230387fb;
// music[5941] = 256'h10fd46fd7d00b80114002b056200d8fe81067903d7fe32feacff27ff6dfd4d01;
// music[5942] = 256'h6c01310b681d2e1c1a19b21dba1c8e1b7b18a411c00eb3128a14ce12eb17ee18;
// music[5943] = 256'h6714de162618ee173a1cb520281cd70a7cfd71fd690099fe5cfbe5fc38ff2d01;
// music[5944] = 256'h4f037f01f2fbdef69bf8f5fb8cfabef715f37af3aef853f99af7fcf479f6b8fb;
// music[5945] = 256'hebf82df440f652f78df555f801fc67f82cf327f5ccf704f5d3f4f4f437f28ef6;
// music[5946] = 256'ha3fbeaf751f0e8eca7f264f7baf1dbeacfeaddeca8ed2deb9ee3aae180e5f2e6;
// music[5947] = 256'h6be920ec6aedb0e615e04ae6fbe868f20206e90313fb69021209fa021cfefcfb;
// music[5948] = 256'h87f429f7bef98af4c6f6f5f287f1d1f2bfead4ed06f03fed3bed2ddbe7c92dca;
// music[5949] = 256'he9c8dcc501c864c7d8c2e5c4d4c4f0be50bffcbea7bdfbc008bfe7bb67c192c1;
// music[5950] = 256'haeb98fbdb4c069bbdabe99bee8bc03c446c24cbef5bde9ba9dbcd8bda4bc14be;
// music[5951] = 256'hbdbd7fc2f5c765c2abc0c7c52fc6f2c58dc57fc503c53ac163c7bad714e2c9e5;
// music[5952] = 256'h43e535e3f5e6cce640df5ae355e849df62de34e50de468e53ee6e9e1caeccbfc;
// music[5953] = 256'h91fc0bfe2701d9fe3c020701b1ff8201f9f9d2f8bafa76f8d2fee30062fd0b02;
// music[5954] = 256'h0306d705ba071902cdf39eeea5eed3ea4de9f4e88fec36f2deef41eb6dee2cf5;
// music[5955] = 256'h38f431f10bf2c0ec78ebd9f3f4f3e8ef3befb0ef30f58ef222eb7df145f40ef1;
// music[5956] = 256'hfff3a9ef5be987ee53f621f6baf20af403f27cee97f01ef25ef736fca4f8eaf5;
// music[5957] = 256'hfaf396f4d1f791edd0e25ce400e305e8fded30e5f9e56de98ae50eebf9e908e4;
// music[5958] = 256'h47e6cae5a4e367e484eed6faacfdfbff70ffb7fd08ff36fc41f8fbf5cff921ff;
// music[5959] = 256'h15fd48fbd9f8c9f62df7d9f697fbf2003603e4fefbecb8e2f0e926ec9ce888ea;
// music[5960] = 256'h17e9d0e672e850e5bce75eeb88e70deb25eb75e87cea18e416e47ee6f6e3abea;
// music[5961] = 256'h1de8b7e18ce95dec18e9b4e751e520e4a4e35ee493e797e743e4a3e68eebe1e7;
// music[5962] = 256'hc2e2e4e58de9aee68ee3bce38be142e21cecdcec85e709edb0eb73e96bf0aaee;
// music[5963] = 256'ha8f08ef1f6eab9ee8beb23e7eae91de312e52cea33ebf6fa5b0205fd85015603;
// music[5964] = 256'hd3fdcef990f584f5c5fbb0ff68fe1afe43fc96f715fb47013103090129fd4303;
// music[5965] = 256'h29feb7e769e3d1ea2aeb89e762ea48ef90e6c6e45ce9d6e7afebc9eb35ec0bea;
// music[5966] = 256'hc1e24fe8a7e96de748eb3deaede857e754e5d8e48fe63dea09e8b8e402e3a7e4;
// music[5967] = 256'h3be728e5f5e673e781e271e25ce377e5c6ef96f600f1eaed6cedeae9b4ece3f1;
// music[5968] = 256'hd3f242f118f3abf761f400ef5fec88ec3ef0d2f2b7f647f52eecb8e963eb7de5;
// music[5969] = 256'h1de2e1f254029cffe502f607640173fe8bfea2ff4c04faffbbfcfd026902a503;
// music[5970] = 256'h9406170074fe20ff81001e079f024af4c4eb8fe948e8bcea9eeebdef83f08bea;
// music[5971] = 256'h67e6a8e7bce5dee99ceaa8e632eba5ed35edc4ec06edcfed45eed0ef96eb20ec;
// music[5972] = 256'hb9f064ee1ef158eeb4e776ed73f2a2f210f03bede2ee2fed01ec9fefc1f16ef4;
// music[5973] = 256'h71f9ecfbccf739efe9eb2eefc4f26efee60c0c0ad405450cde0aed07ab0c1e0d;
// music[5974] = 256'he5081505a905110b6c0bac0577ffd001a21436228f1df21c8c1d9d1592180e1e;
// music[5975] = 256'h371832173e1a9f1c371ca6169d1a341d4b17b718fa1ac31d6d1d250f8b026a00;
// music[5976] = 256'h7301b5000801f60071feb8002f0299029a04aa008ffd02fe49fe8bfe49023006;
// music[5977] = 256'hc2ff8afe350475022e020304a20670072d03a8011d018203100204fabbfc4d04;
// music[5978] = 256'h8804d2039804a1ffe3fa1effa9022c08b10970049708f709cd090b0971fdaaf9;
// music[5979] = 256'h5df553efa6f327f191efbbf6f3f98af3ccefacf449f158f29bf304eae3f68108;
// music[5980] = 256'haa0aa30953012900b102ffff44037205e0039a00e003b409e9034b015502f502;
// music[5981] = 256'h8c06ef006a008a0546f8acebececc1ed96f086f038e951eba6f2dfef47eb3dea;
// music[5982] = 256'h52e6b1e628ee66ef05ec30eb05eda6ef00eabee5f5ed62f077eb0dee79ef78ea;
// music[5983] = 256'hf1e9a2ec9def5af0faed27f143f0daeb92edf4ec1df070f0e3ea38ee7aef39ef;
// music[5984] = 256'heaf08ef2a1f4f3f090f3f4f618f5e1f709f3b0ef36f35bf128f0c9ee44eee2f1;
// music[5985] = 256'h77f1caf1b9f740f7b4f73a094312aa0a7907cc036e01eb046702c9fee2010404;
// music[5986] = 256'h1c05ce064d00cbffe00897063104020a000ca508c7fcb3efd4f04cfbbafe6bfb;
// music[5987] = 256'hf5f8aff961faddf6fbf852fac4f4c9f8abfc29fcbcfe8d0094059108ba08bb0a;
// music[5988] = 256'h020e0d10db0cf70fbc156f15b812a20b960bce0c96087e0d5a145c0f73030b05;
// music[5989] = 256'h9f0d2b0c0711a915e616db1bdb153c12301477120215870ead034902bb008ffd;
// music[5990] = 256'h54fadffb4cfe13fa6cfa56fbf2f993fb94f7baf2adf53306ca18b314200f9215;
// music[5991] = 256'h5f161518db1cad214828d2284927182aea2b322b222da22f122f312fe335b03c;
// music[5992] = 256'h5232502349201a1ffd216424412435299528a327272a06285027fe298d2d042b;
// music[5993] = 256'h4a29e82d172a67274b2a31272028ad2c3d2cc12c0c2ee229f727302d8f2d202c;
// music[5994] = 256'h6f2f532def29d62b772b042cf02f682ec02a0f2d7f30c92f5130c43537391837;
// music[5995] = 256'hf4333937d2410646774123403641274279443543cf3e733ee53e4a3b8c3c2140;
// music[5996] = 256'hed3b3f40f74e7e4f454a5d4b2649ab4a4a4d194b334e204de048aa4c954b1246;
// music[5997] = 256'h954681481e48cb469a46f7485447bc39fe2cc72d802f382b81285b29732aca29;
// music[5998] = 256'h9f276e26542684252d268b268526a828bb2546215d21f922df255d268624dc1f;
// music[5999] = 256'hef1b701f6a1eb11b001e8b1baf1a9c1dd01bde19bb1a501a3818ff1630188019;
// music[6000] = 256'hb516b619aa20911d7a1e2221f01cc61e90180e0b30095b0a180a38091b071905;
// music[6001] = 256'h9a0543088105d102d7035d031c022e036a0d0c16ae158115c8140017cf181818;
// music[6002] = 256'ha31a01176515161afd17291596142316181a0a1c5e1b6c182f19e312f101ebfe;
// music[6003] = 256'hc8036302f50016012703db0282ff23fefcfdc3fe24014f047401f0fdb8029903;
// music[6004] = 256'ha4002f028d031c03db00ffff2600cafdc4feec005bfec0fc430033033100fffc;
// music[6005] = 256'ha7fd35fc7ef95afa2afc5efb6cfa88fe8d02d2015e01a1001e0409088f02bf00;
// music[6006] = 256'hee0003005105a702b9fe3c019c017f032a022302ee04ff03e102cefc0004fe13;
// music[6007] = 256'h16119211aa162e12571364162d13720fdb10c7127f132316f1134f13e7151e17;
// music[6008] = 256'h7c188116071b9419c505c2fcedff2700cefdeffc0bff84fd48feffffdefd80ff;
// music[6009] = 256'h43fcccf7fbfc840149fe5cfacdfbc4f9faf5fdf668f648f86df9bbf583f574f6;
// music[6010] = 256'h88f5f7f278f33bf68bf2d0f152f732f6fbf1cbf1d2f1faf3e2f614f3d3f3daf9;
// music[6011] = 256'hbef60ff205f67efef9fdd0f51cf464ef39e90be9c0e5f6e32de4a6e61beb13e8;
// music[6012] = 256'h97e6c6e8f3e7e5e490e59df51902ecfd2bfdfcfc61f8f9f668f632f90bfbc8f6;
// music[6013] = 256'h4ff61cf64bf15bf135f0f0ebf0edc0ed9ded7befd7e006cfb2cd11cd20c9b7cb;
// music[6014] = 256'h82cbf7c5fcc687c90bc7acc579c305c1d3c247c3c8c1dac25bc362c182bf2abd;
// music[6015] = 256'h46bd1ac13fc02dbcf4baa9bcfec15ac2cfbe0bc208c4f3c295c4ffc3afc4c8c7;
// music[6016] = 256'hfac465c28cc665c962c950ca28cc20cdaecbfbceddd1a9cfacda62e695e200e2;
// music[6017] = 256'h9ee497e362e281e353e5b4e2e5e1cadf7edf01e5c8e1efe9ddf9f3f62df78afb;
// music[6018] = 256'h2efa25fc5afcb8fb2cfcb4fc0efb37fb150002fdecfa8d0044035a025dfe85ff;
// music[6019] = 256'h37fe38f0e3e7abe9efebbfeb2eec05ed2bec7fef3ff11cee52ec24ebf1edc9ef;
// music[6020] = 256'h3eee84efafee27eff1f3dbf221f130f58df55cf2bdf108f1a4ef89eeaeefa4f0;
// music[6021] = 256'h0cee08f066f400f3ecf1e7f15df10ef330f30df424f807f8cdf9a5fc98f8b7f9;
// music[6022] = 256'h86fbc8fa73fdebf231e723e8f2e70fe96cea9eea09ea7de79fe91ae750e562ea;
// music[6023] = 256'h77e7d5ea73f8cdfc47fd3bfe42fcb7fa77f8a6f9d2fe87fddffb61feb7fb58f9;
// music[6024] = 256'h93fb5cff71027700d6fe8400dcfe68f3eee535e75fea30e62ee836e9a8e5aee5;
// music[6025] = 256'hfee626e8e5e50be5f5e9aee81fe618ea72e93ae7bae679e32be5f9e886e88be8;
// music[6026] = 256'hb3e7ede6e4e6bae341e3a0e755e75be45de412e222e24ce4f0e14ee618ea7ee6;
// music[6027] = 256'h44e9d9e80fe43be756ebbeec2bed5dec44ebc8eb96ecd7eb65ed01edceebdfed;
// music[6028] = 256'h7beefbed09e980e576e9a8e807e4bae6b6f487000802ff01d1ff0b01be002dfb;
// music[6029] = 256'h6bff1100f2fc96ff98ff42022401bafdddff59001b016e0099020afd2be91fe6;
// music[6030] = 256'hb3ea05e716e7f9e4d7e38be5c4e34ce518e939ea1be961e7dfe507e8dceb23eb;
// music[6031] = 256'hb2eba1ec0deaf7e837e5a4e332e904ea34e92fec1aec5deca4eb79e6c3e6caea;
// music[6032] = 256'h41ea69e7f6e6a3eae2ec7fec03ed04ee21ef2dee18ec8beb00ee7ff1a7f04ff2;
// music[6033] = 256'h7af5f1f1f4f022f2b2ee81eff8f399efbae922eec5f05cee7becdbe8a8f2c705;
// music[6034] = 256'h53073403c605ab04bf053506b1fff8fec802c9032203f7007201d703fb03b803;
// music[6035] = 256'h02069706c50493026ef580eb00f023ecd4e9e8eca5e8fbe9cdeb52ec09efa3ec;
// music[6036] = 256'h9ced7beeb2ecefeb87eb13ef41ec7be8bded8fec23e91febd4e9b1e908ee10ee;
// music[6037] = 256'h19ed96efdeed86ecbeef82eeb7edf6f1f8f130ee41ed68ee02f1d7f1d7eff4f0;
// music[6038] = 256'he1f280f3c6f30cf6adfb1ef9a8f8d106880f9a0e9a0b450887064904a0068e0a;
// music[6039] = 256'hb908f705e8057906fa073714d4219b21bb1e8d1d0e1c151ba9179518f71b3c19;
// music[6040] = 256'h4618461df11b7318891bbb1be61c931d3d1acc1d7916d3050e03650313025200;
// music[6041] = 256'h4b0020053102effed500b7ff7c02b00366002f03a60532031f032d0544068d07;
// music[6042] = 256'h070687026b043d058f01cf006cff67ffc00343054004bd00f5fe5f02ca0068fd;
// music[6043] = 256'h7f00ea0211016403f006b00294006a001000f4051a06b707f7091cfc62f5a5f6;
// music[6044] = 256'hbdf34ef649f47ef0c6f0aeeefbf0d1f125f038f01bede8f73f0c3d0b92043e08;
// music[6045] = 256'h8d06ba020b024501ac012d030e06f004120563076704d70559096c097108bf05;
// music[6046] = 256'h7c030af7edead7ecceedfbec5bedc4ef02f184ed49ef65ee8cebd0ed9febd8e9;
// music[6047] = 256'h1cea73ec97f0d5ed25ecaceee3ee5fed3dec26ef4af0c2ecf1ecb3ed1decc3eb;
// music[6048] = 256'h1ce97ce933ee51ef78f1dbf0feec1def4cef2fee84f110f42af1a3ec43ef62f2;
// music[6049] = 256'haff092ef39f13cf5e6f5dff609f761f4c2f5c2f6e3f390ebd7eac8f3e6f00ef2;
// music[6050] = 256'h15f680f70c0a3c124a0c521051107e093a047c03b702f3ff8800aaff5c010704;
// music[6051] = 256'h4b020104b3064507b904a604e80872ff3bf1a1eeb3eeddf368fce5fceffaf7f8;
// music[6052] = 256'h35f682f7f7f775f616faf5fffc01e202e40401048f05eb09310ad40e2f12460f;
// music[6053] = 256'h59127f11f60d6d128313cc107c0fb611ba15261566155f0f2f02ef010b08b50b;
// music[6054] = 256'h751190126712cd15ed1431107c0dc40bf4076d04ba0268034d04a9fe28f864f8;
// music[6055] = 256'h5afc48fcb0f8e1fc35ff84fb96fbd2fa3d08761a9218e618451c511b8720e320;
// music[6056] = 256'hd81d351cf51c6a24e326bc2493266928c52ae22fb5319e315437f2336123411d;
// music[6057] = 256'h49216423402474243d247a243528bd2a23277c26d729ac2ce22e892c9f291b2b;
// music[6058] = 256'h002d482ddb2dc83004307a2dfa3000316e307932902e872cc82cff2f2934052f;
// music[6059] = 256'h422fbe31422d4b2e752fa231a03514329c2f8530da2fd52ffd2fc52e3c2d092c;
// music[6060] = 256'heb2fb83d4845ba416b413841414021409f403a44f0413a3f6e3f5b3cbd44c954;
// music[6061] = 256'h89593d58dd5667543552a3518d51d74d204c394f774df24c5f4e444939473b48;
// music[6062] = 256'hb14793468b468e49953ed72f432fb62c962c712d31295f2bc4296027462bee2b;
// music[6063] = 256'h102cf9292a26b026c6271e25ac23fb267b26ed251829a5264f24f422bd1e871e;
// music[6064] = 256'h3d201a20611f7e1ef820ba22101e651a921c471ff91b6e16ac18ba1a971ac81c;
// music[6065] = 256'hb41be11c8a1c401bae1d291a8e1d0b1a1207fb058509df069a08b9079a07b306;
// music[6066] = 256'hc0073308870541068e04f60ff31e3c1c4f1cbb1c1c1ce81e9a1b241bec19eb15;
// music[6067] = 256'hc11596163a17c416c0186e17ba15541a2918ce173315600465fd770086fe64ff;
// music[6068] = 256'h8b03c901f8fdd001ec0371ff9bfe2fff5efe7cfffe011603e400d6ff8d01f101;
// music[6069] = 256'h6a000bff69ffc4fee4fc93fe6efe2bfbb0fe1a01d5fcb6fddbfe24fceafeeeff;
// music[6070] = 256'hbafb3bffb404ba014301b403f700080067014301e500ee00e702ee0099fd8200;
// music[6071] = 256'h7e03d8047c0343018a0206028e035a05f60146ff0cfd5104ac140f1bf919f61b;
// music[6072] = 256'h9d1e021a1116ce1aa61934169d142b1051137b169615da1518148216a317a019;
// music[6073] = 256'hb01bf50ae8fcd1000a03fd00d1fda5fb29feec010402e0ffe3fecdfce3fd66fe;
// music[6074] = 256'h3cfc7b00ebfe10faf5fc60fa24f6c9f36ff3bef8f4f591f312f958f76cf739fb;
// music[6075] = 256'ha4f869f9a8faeaf6bcf665f627f51df5e5f26cf420f485f1f9f4a0f236ec5ceb;
// music[6076] = 256'h07ef83f471f019ea80e92ae860e873e783e864ecc8ebd4eca3eeb3ef67f093ec;
// music[6077] = 256'h58e7b5e849f846067a0635062405580374039200e2fd55fd48fdb0f8ccf4f8f6;
// music[6078] = 256'h64f62cf54ef401f236eea1ea97ef31e779d058cd6cd157ced8cdf0cce3cae5c8;
// music[6079] = 256'hb3c81cc94dc685c48dc58cc6edc576c59cc325bfe9bd6fbfecbfb4bd4abc2fc0;
// music[6080] = 256'h0dc2b0c1f4c290c39fc57fc4a3bf30c1e6c498c305c38cc516c54cc105c1c2c4;
// music[6081] = 256'h77c57fc5bac9f5ca48c843ca07ce69cb85c8a1cabcc8acccc3dc30e46ce342e5;
// music[6082] = 256'h59e887e84ee37be2f1e32ae52de7d1e286ea3ffae9fb17fdc7fe0f0074038300;
// music[6083] = 256'h8b00bb004dfec201fd0240ffacfa85fc23036701cbfecdffcc005c0047f534ea;
// music[6084] = 256'h67ebddec13ecb4edb3ede2ec17ed0aed52ef12f0efed0aef98eeb6edcdeeb7ec;
// music[6085] = 256'h86eec6f0c2ed21f030f323f1e9f002f24bf264f494f45bf0d3f114f5cdf0a5ef;
// music[6086] = 256'h92f151f1fff1c3f2d7f376f34af527f802f73cf99ff8b2f416f750f647f382f3;
// music[6087] = 256'h2cf513f603ee89e648e925e9dee66ee992eb72ed0beee1ec57edbbe887eab6f9;
// music[6088] = 256'h24ffb1febf0102027304a804260422048bfdcffabdfebb01b1fd49f992fe7700;
// music[6089] = 256'h65005e01bdfd98ffc1f74ae57ee32ae77de525e73ce919ea17e8a5e4a3e5ebe4;
// music[6090] = 256'h3de288e6eae857e53ce74dead8e7aee60ce64fe448e8a8ea84e58be597e898e9;
// music[6091] = 256'hadea46e61fe398e459e5f0e628e6b4e4d4e247e267e63fe636e723eabee616e7;
// music[6092] = 256'he2e848e639e622e8ebe74ee65ae645e64ee9e8ecc6e8eee81cec4dea13ebcaea;
// music[6093] = 256'hc3ebc2ed89eb20eab7e9c1f42d04f00235ff6503ae05a30155011405c0fee2fc;
// music[6094] = 256'h68001efe4602bd03c1ff0700420072008ffe7c026c02e4f0ffe600e817e627e4;
// music[6095] = 256'h37e3d9e3f8e31ce572e810eba6e95ae42ee4d1e781e95ce9b4e90aea50e796e9;
// music[6096] = 256'h81ebfee846ebe6eab5ecdeefcaede8ee27ebe7e8ecec58e90fe816e94fe7cce9;
// music[6097] = 256'h5aecc0eb97e9d6e7a9e92eec24ecf9eb74ebb3e9a9ebeeed67ecf2e84ce8e5eb;
// music[6098] = 256'hceea61ea27ee6eec1cecdef0edf3d0f125f22ef576f06ef486010106b007b706;
// music[6099] = 256'hab06e3065b044f0713073506e8065d047c06090555036706b803df03c9055e07;
// music[6100] = 256'h410870f8f9e676e7f4eac9e9e9e875e830ea50ee30eeb2ea1cec9eee13ecebe8;
// music[6101] = 256'h2dea58eee7ecbde97cec99ea28e890eca1ecb5eb7cec31ec1eee92eb4ae906ed;
// music[6102] = 256'h1fec86eb0eefebec0de943ea41ed2bee2ceda5ecfaea27eb59ef07f188f12df1;
// music[6103] = 256'h89f09af211f0deeff2f4d8f9a504a709a606680a490ccc066f06b00c9e0c6c0c;
// music[6104] = 256'h2b0d8e08b614f922d51ec31f6c21c31fac1f781c411e271e5c1cc01e241c471a;
// music[6105] = 256'hcd1c141d391a301a841b6d198c1cc6168904e10266055effbc02f70471008d00;
// music[6106] = 256'h3a001c009502bc0320051c045103e70395026c040f06c7059e04030185031706;
// music[6107] = 256'h3a032f0306036702cf054d07a802550126034cffceff3303dc02670284ffab01;
// music[6108] = 256'haa039afe990004049601c20092035804ecff47fffb027805b5fff5f089ec85ef;
// music[6109] = 256'h28f0b6f339f2e7efd0f1b8f141f19cef6ef9760ae80a8c09d40b8707a3063206;
// music[6110] = 256'h3d0619083c07a00ab50a59071a098509bb0a8b0b5709d905490376046cfa71ec;
// music[6111] = 256'h7ceca1eb18ea89efe4ef4aeb8dea15ed1befbbeeebeb26ed8aefcaed75ee7cee;
// music[6112] = 256'h3ced48edcbe927e951ed7ef0e6eec0eb48eca7eb41eb69ec58edd7ee6dede7ec;
// music[6113] = 256'h33ebd6e976ec0eeb4fec27eec7ea70ede8efd2ebdfeac5eeb5ee06edd6ee9fed;
// music[6114] = 256'h7cf021f5a2f146f1f2f294f1aef2f8f368ef9ae8fceaafef10f1e1f2f5f7c307;
// music[6115] = 256'hb810fc0b6a0de60e750cb50942060f09380b990654058209720ace06a2055d08;
// music[6116] = 256'h980b8d0a3f09a60b930385f459f248f357f115fac900cdfaf0f851fa86f529f2;
// music[6117] = 256'h1af5c3f834f8bdf7a3fbc800150411052408d60da4102b11a111fd1212157a12;
// music[6118] = 256'hbb0e2d103011c711d212930f2b0d2f11ec16940d1dfe7c035e0874053c0e7b11;
// music[6119] = 256'h441177163a14f30ff10cbf0b950bf007ff0463fffefa0dfd8efadcf55ff61af8;
// music[6120] = 256'h7ef70af53df672f9defa3806d114c3165e17a0173e155c191f1bfc19be1da521;
// music[6121] = 256'h1e2223247b29122bda2e8732bd2eed320837e1341534242a48206d1e701f6b24;
// music[6122] = 256'h49258c24b32681270b2849294b2a1a2a9a2b3c2c962a402ae3282d2ae22af129;
// music[6123] = 256'hb12efa2fd92e902f092dba2dd43053305030e030612d922ba02e982de12d5230;
// music[6124] = 256'h9a2e5f307c311c307730132d71298f28ea2b5e2e832a9d2c8731653252320b2e;
// music[6125] = 256'h2c3276400043173e6e3fce40c8406b425641b63e413d02422d5013590b576f53;
// music[6126] = 256'h545001503752e550294dfa4df64e604d544fef4ec64dc14e294cb54dda4c5349;
// music[6127] = 256'hd049c93b202c162ccc2b832ace29ff28ed29f9273f28272c9b2ba227cd26f426;
// music[6128] = 256'h162622268e24cd25d427c425a828332adc260b26e82445249a222d22b0235120;
// music[6129] = 256'h6921a123a21e181db31d191db81d771c181a5f1a071dfc1b8d19331a24183a18;
// music[6130] = 256'hef1ba11b561f3a23251d6a1b561a660e71076107c70549050e0647072e05d205;
// music[6131] = 256'h7d08dc05b00fb71dc21d9a1d451afc16b71ab918e219fe1ebe1bc81b911fe61b;
// music[6132] = 256'hb41a101fc11cf61abe1def1cfe1d2d192609bb000301560045006900a2feaafd;
// music[6133] = 256'hb7ffff00be007f00dffe39fdd8fcdefb3efcc7ffe1fe4cfaa7fb4ffdb7fdf800;
// music[6134] = 256'h5a01840099ff52fc89fb89fc43fdd7fd6dfce8fb82fd33fed1fe26feb3fb0cfc;
// music[6135] = 256'hbbfd7afefafd70fb3bfb7ffca5fd7e007a025b036e024602c6035b026a019f00;
// music[6136] = 256'h42010a03dfff1501f7016efe4501edff12034914571ca31b7219e916ba195a19;
// music[6137] = 256'h24170717c415fc16ef16c4155816ec156a16f416e4174a17a8160c19b50fedff;
// music[6138] = 256'hcdfce5fe0e00b600faff7c00f9ffcffd7ffb9dfa00fc09fb73f828fa0ffe36fe;
// music[6139] = 256'h65fc06fb21f834f6d9f53ff5caf43af428f5c2f556f51bf608f50cf5f2f622f5;
// music[6140] = 256'h7cf332f3aff19df110f2d4f146f143ef8bed41eddfec5cebd1e8c6ea83f418fa;
// music[6141] = 256'hdbf4eaefb4edbbe914e72ce50ce5f6e6c1e5f5e615e95ae661e704e7dee793f8;
// music[6142] = 256'hdb05b905d204b6021902b50005fefcff07fff8fc7bfcadf9a7f841f8f7f751f6;
// music[6143] = 256'hb4f392f3a6f2e9f2bfea7ad9e6d214d0f0cbe8ccaccb8eca23cb7fc959c8b1c7;
// music[6144] = 256'hdbc527c4f4c31ac30dc1f9bf34c0a1c009c077c1b0c1aebe23bff5bf4ebfffbf;
// music[6145] = 256'hdebfc8be8fbd95bd09bd6dbdd4bfc1bdbdbb28be5bc19dc2d6c07dc087bf70be;
// music[6146] = 256'hedc044c1a7c3e2c67fc53ac7cdc75fc62fc969c799c812d642de17dff0e01de0;
// music[6147] = 256'h8ee1d6e24ce1fee280e281e988f921fd13fcc1fe14fe9efdf4fd87fe0dffbfff;
// music[6148] = 256'h61014901f1011c026c02d5042104c203b70362040d05e0f801ed7ced1aec43eb;
// music[6149] = 256'hfeec36ed27ef4def98ef82f08bee7deebfeebdedfbed86ee95f01ef25bf2f7f3;
// music[6150] = 256'h05f49df240f204f29ef38ff4a6f2aaf257f36df336f399f0d2f079f287f2bcf4;
// music[6151] = 256'hb8f46ef299f218f4a5f3f2f0b8f165f36df31ef50bf6b5f53bf583f834fbc6f8;
// music[6152] = 256'h57faedf581e9bee6cee608e408e4b9e481e594e735e6e9e652f5cbfee6fa53fd;
// music[6153] = 256'h9a018d02c10179fea2fdccfd7c00e70035ff7002e501e9018902f5ff5f013402;
// music[6154] = 256'h280451fddeebb3e801ea49e6cce6e8e6b4e7d3e7b8e6b4e755e73be782e7c8e7;
// music[6155] = 256'h24e8fce52ee647e7f8e496e6baeac1e91de9d7e861e5c9e58ae6c6e351e421e5;
// music[6156] = 256'h90e486e5dee633e87de764e633e631e540e514e5d3e39ce2dfe2ede5e5e556e3;
// music[6157] = 256'h3ce33fe340e34ce3e4e41be881e82ce992e9e1e712e9a8e9e5e842eab8e9c7e8;
// music[6158] = 256'h98e7f3e60bf1edfc8efe45008703f00432067c04d902700166007d013c01d802;
// music[6159] = 256'h25048c033104300233012e012502f40006f2c0e637eadbeb28ea9ee8abe71fe7;
// music[6160] = 256'h32e6d8e6dfe681e696e6fce53ee7a5e84ae784e61de80ce910eb91ed10ecbce9;
// music[6161] = 256'h09ea0bebd7e9a1e92aeb08e9c4e8afea71e9b2e77be61ee8d7e837e7c3e741e8;
// music[6162] = 256'h21e900e812e7f6e83de719e7e9e85fe9c9e99de8c7e848e9b4ea95ec17ec3ded;
// music[6163] = 256'hb8ec77eb39eb42ece2ed0feb8aecefebf6ea3efc4206cf0294056606d0062608;
// music[6164] = 256'h8c07c00711066c061007610626080009d607cf055e0616078d07a409f7fe17ef;
// music[6165] = 256'h0eee61f065ee9ceddeed3fee9eecbaea89eba6ecceebe2e926e964e99dea95eb;
// music[6166] = 256'h1eea37ea08ece9eba8eb9ceb62eccdecd5eaeaea8feac1e83cebf2eb8fe9dbe9;
// music[6167] = 256'h73eb52ed74ec9aea9beb3aecb6ec0dec79ecb3ef80efdeef14f128f004f02eee;
// music[6168] = 256'h13eeb8ee2eee91f14bf346f89502b203ba0009040807ca05c606bd04f800a40e;
// music[6169] = 256'hb11c611bd61ce91d171ed021dc200d20611fc21c291cc21c061e2f1dcf1c911d;
// music[6170] = 256'h581edf1ef01bce1ea21dec0bfd017d03e903e604170462042a040b025e04f904;
// music[6171] = 256'h170365045004b401bd0070029d0337023802ee04ac04ed02e703b80331034403;
// music[6172] = 256'hd901c30003ff4eff9c0047ff3e000f00edfece000a0092ff03028603a50277ff;
// music[6173] = 256'h5ffdb3fc9ffdacfe96fe5b00bd0064009101c700e902440411fabdf0bdf249f3;
// music[6174] = 256'hb4f025f01aef73ee13edc7f45a057109a407fb07bd078e0b5c0c970bdd0b530b;
// music[6175] = 256'h940c00096f063209d90a920a1e08b8091d09b2070a0ba8fe7defc4f0c0f1a8f1;
// music[6176] = 256'hedf19fee98edfeeeb0ee0aedf8ed47efb7eec6ee91ed0aec74ec75ed91ecfceb;
// music[6177] = 256'hcbee25ef9ded8eed27ec79ecdcec16ea69e9f6eb84ed67ec69ec59ed91eca5ed;
// music[6178] = 256'h36eea8ecbcee06f1fcef3aee93eb93eac2eb2aeb2aeabceab3ec61ee0ced9aeb;
// music[6179] = 256'h48ec3aed9deeadf09cf45bf7ebf102ea89e99dee7ef128f50504b911f3110f12;
// music[6180] = 256'hef12a6102110c40eb60ea90ed70b450b0209a9068b087908a80728091109a309;
// music[6181] = 256'hf60cc006dcf7d6f3dff534f207f4bafcd5fd13f9fef8d9f81ef68ef529f51bf6;
// music[6182] = 256'h28f909fc81ff32022d044206290a350e5a0ebc0fbc111010ca0f4110db0fda10;
// music[6183] = 256'hed100e1053104a10f80f6b133816530ce4013c072d0c3c0ce8108d111e118312;
// music[6184] = 256'h1c10a10fdd0d100920056f00fafdb6faf2f634f793f721f8e6f78bf571f376f4;
// music[6185] = 256'hd5f66ff699fede0dd6125212c71344161f19121c941f1e211f23cd24ba25aa29;
// music[6186] = 256'hd629d629f92c992df72f41311533ba340e29a81e1521c0221b232224f222b423;
// music[6187] = 256'h0027d627c42669270829952ab42a352a912b8b2b762b5d2c9f2bf92ca02e602e;
// music[6188] = 256'hfb2e9e2e222eec2d072d1d2d2d2d1d2de02c002cd42b082c442c752da72ec72d;
// music[6189] = 256'h092c392bea29732728265327d22794283d2a3a293229e82999298e2a6e281f2a;
// music[6190] = 256'h3735373c183b8439e23832395c3ba5390b3b184af6527f503f51db4f714e6d50;
// music[6191] = 256'h76500650664f774f424eda4ca34d7e4b9f49ec481248b24719468b46303f1930;
// music[6192] = 256'hfa2cbf2e8a2ce62c932c752ab0296f290229a32840286b272727ad26c025cf25;
// music[6193] = 256'h6225e024ab24c1233a241b25e923f322fe22752277214b20b51fb01ff61e321e;
// music[6194] = 256'hfd1d741d9d1df91e8a1e291d5d1db61ce11b991be01968191a1a201acb19ea18;
// music[6195] = 256'h121861172f18fc17f416eb17f3101306730355048f0690064505eb052c05e10e;
// music[6196] = 256'hbd1c411df11bbe1c0c1c111d461e441f181f0b1f2e1f6d1eb81e681e921e041d;
// music[6197] = 256'hfa1a511c171be11bd41abb0cc702b403310389020303890141003500f8ff2a00;
// music[6198] = 256'h7200650088012c02a8017501dd006c0021007fff8cffc400d701880100018801;
// music[6199] = 256'h4d02af01ce00e7005700e9ff78ff25ff7300a100c4ff74fff9fe85fe10feb3fe;
// music[6200] = 256'h45fe66fc79fcdbfce1fc49fde3fd8afe90fe06ffd2fed3fe53ffc7fd16fde8fc;
// music[6201] = 256'hf0fd4001840295039d027d050314d01a5f17d017cc17ff19681ea01df61bcb1a;
// music[6202] = 256'hae1983192b19eb184119141ae118a41744179617e81929126904d502a104b803;
// music[6203] = 256'h8c04d102eeff10ff05ff0effbefe96fef2fd80fb89f8c4f988fd19fd98fa71f9;
// music[6204] = 256'h75f8caf7d1f723f8d5f6daf404f540f58ff5c4f6b9f670f674f661f7e6f818f8;
// music[6205] = 256'hedf67cf6b0f548f5dcf447f42af336f261f009ed7aea3aea67f0b4f40befbbeb;
// music[6206] = 256'hd5e928e556e349e075df16e228e275e37ae531e888e965e913f51902fb01a301;
// music[6207] = 256'h5402a10045017c01cb003400a4fff8fed4fdccfd56fc88fa16f92bf7a7f54ef2;
// music[6208] = 256'h84f2b4ee51de72d577d5e6d214d22dd1bece2acd86cc06ccf5ca61ca25c9e6c7;
// music[6209] = 256'hfdc6cbc551c570c4eac3edc2dbc1b4c1a4c00ec114c2a0c12dc1a0c0f4c0e5c0;
// music[6210] = 256'h67c008c00ec0a0c145c14ac0a3c022c064c0d1bf70bf91c008c092c039c101c0;
// music[6211] = 256'h30c0cbc078c122c265c270c308c4a8c5c3c57fc44dce4cda84da3bdbe9dc97dd;
// music[6212] = 256'hf1e2b1e261e60cf69ffb63f99bfaf3f940faa2fc55fd8afdb6fe91ff82ff3200;
// music[6213] = 256'h42003d01e90273025f0379020b01df0177f894ec23ec17ed21ed88ee70edf3ec;
// music[6214] = 256'hb2ed0dee65ee16ee47ee7eee4feefeee3eefaaee84eeceeec5ee06ef08f026f0;
// music[6215] = 256'he2f0fff231f320f3f5f3a2f352f3b7f30ff5e1f560f4cef336f43ef487f4ccf3;
// music[6216] = 256'hc1f33df45ef438f531f5aff5e0f426f3d8f4c2f5faf543f616f61ff6eaf2f2f3;
// music[6217] = 256'h7bf3b1e80ce40ee66fe62be628e579e57ae7d3f2affed9fd00fea0fe8dfde2ff;
// music[6218] = 256'hc4ff8b001c024f02c502020240029401cf0108038e02d702b10170012ffc30ee;
// music[6219] = 256'h4ee99bebf4ea18eb76eae8e8d2e85ae9c6e992e90eeaaeea87ea98ea61ea14ea;
// music[6220] = 256'he0ea45ea9ce81ee97ee979ea34ecebea44ebb0ecdaea64eab6e9dde822eb5aea;
// music[6221] = 256'hf9e75de8efe7d5e604e644e625e7bae611e744e7ffe6e8e6f1e5e3e5bbe4a4e3;
// music[6222] = 256'h87e5efe542e55ee4d8e3aee53be698e683e77de7b0e85de89ae96eebbde8fff0;
// music[6223] = 256'ha3ffb9004d0042027a01060411049802ab032c0350034f032003c3022702c302;
// music[6224] = 256'haf02ac03a0020003360383f409e90feb8cea69eb9ceb12e8aae872e98fe8c4e8;
// music[6225] = 256'h76e9f8e9c5e943e96ee8f0e750e765e600e7c0e855e971e908ea98e9fce959ec;
// music[6226] = 256'h1eee76eecced09eeededf0ec0eed32ed66ed3bed6fece0eb57eb01ec91ec9fec;
// music[6227] = 256'h99ecf1ebfeea42ea18eaffe721e784e8b3e689e612e771e6d5e89ee9fce95bea;
// music[6228] = 256'hcbe912eb02eb5fec60eb48ec2afc2a06c1039904e404eb069408570683077107;
// music[6229] = 256'h27076c08fd07cd0848089d072607c60675079f060109b80236f157ec31ee5eed;
// music[6230] = 256'h14ee35ec76ebdeec63ec7aec58ed0eedebec56ee58ee35eed9ed46ec86ed0cee;
// music[6231] = 256'h4bed37ee5bed8bedaaeee8edc4effff12af2a1f3d2f26ef129f222f007ef70ef;
// music[6232] = 256'hf4eee3ef51ef8eee51ee75eed8eec6edb9ee52eeb7ed51eee8eb0deb55e9aee9;
// music[6233] = 256'hbaec39ecc1ed0ded09f1cbfe4a041a03cf03990478035c031d05d40489070906;
// music[6234] = 256'hf5069119ef2416221c230e244b23cb23412306239a239121861fd51ecb20ca26;
// music[6235] = 256'h682861273a272f254125fd22f61fe71b6d11d80ac708b809de0d060b21061503;
// music[6236] = 256'h24ffb3027a0b260d3f05e1f63eeec6f25ff91af7fceb31eb04fe500d4a10380c;
// music[6237] = 256'ha70bef1684194e0a36fd2f01fd098f0057e68ec89ac1fbdd73fc7409ce0cce0b;
// music[6238] = 256'h670a5909dc076803acfe5500f6036d055a0df216f21220084e048b0e2d1f6921;
// music[6239] = 256'heb13e507170d621dd926131f0d0478eccfe530f1720ff62b5544f44f3c3c4623;
// music[6240] = 256'h7b1aca25e93ebc4c7243842c981b3f17f6162f18d41a0b1be317bd1c71295c30;
// music[6241] = 256'hac2a01226d21d613aef916ef07ea0ceca1011815dd16c80ba5fbb9eee5e71ce9;
// music[6242] = 256'h9ef6f1048c0b8e15d318880c07fb6be80ce228eddbfeef10cc1da92ab8362232;
// music[6243] = 256'h91233922733198453c4ed83f78290f1bbf0e06fd80e71ad584bf5eaa5aabf9b1;
// music[6244] = 256'h4da59e9c4bb084cac7ce54c544bddfb99fbd51c014be0bc533d966e91ded23f2;
// music[6245] = 256'h58fd5f05f2115627e0335c32592d563ab55fa375f86fb2697e692475b479de60;
// music[6246] = 256'he2535f604a5d6e4d154dd955a7574d5bb16188546f3c163ade53ed6ce35b392e;
// music[6247] = 256'hdf1dff2c8b35063bca523466f35609377c26322bfe3474362b358c366b39013e;
// music[6248] = 256'h53454752e061ad6dac753e7617657246a02cb01f981ae510bbfd81f232015f28;
// music[6249] = 256'h5a4a16425029e02e583261164dfe34037c21ef351828b412d2118b2b3a3a0c2a;
// music[6250] = 256'h9c25252e6731562f72277528fd2c852662168a112e260c2d051da61c672fbc30;
// music[6251] = 256'ha31879104c1eae326247b7477142be433e423442ae397e20450474fa3f043b0e;
// music[6252] = 256'hc611751326202735e938ae20e7fa6ddc30de0c03c512690124f472d3b8a85099;
// music[6253] = 256'h249bb1b3d8d519d936bde3a4b4a817c2c0da62e4deea71f53102e4111a0fb2fd;
// music[6254] = 256'habee00dfafdb20e340db56be67a4cd9f06aaf5c0f3d975e0a3d79fd3d1d3a2ce;
// music[6255] = 256'h90d051db33dd40c973ae46b056c172d009f04114b8210b12caf13ee1b2f7cf1c;
// music[6256] = 256'hfc2ce72d87284824ee2990323b3fd7478b447a447d48dd4aee49b235b2151216;
// music[6257] = 256'h4932f244194d924d6a553d6d23791474ae5f653a87215b2da24be05a6156bf44;
// music[6258] = 256'h7736343e833c1f24102191314833aa2fe72e132a14296a26d91ec51d9422ad26;
// music[6259] = 256'hb521a9167a0ef90f8b1b861489fb8df01ef178f55bfc04084f1a381aaa0299f0;
// music[6260] = 256'h3df006f97501760145f659ec37ea54eb8cecf9e56fe2abe896efe202eb10d903;
// music[6261] = 256'h7bfa3207a7179c1427054df9f7ed0ef84d168922171941112d1b7729a022cb07;
// music[6262] = 256'h5bfbb213bc2b2228501a2215c020ec3149337121db1fe52f462ab724e2286421;
// music[6263] = 256'hbc241f3fd15a7e57c835c810c5f8a6fae10942165322b7345749fe492f46884e;
// music[6264] = 256'hba53544a2834d72ab22bf82d6632f91283e45bd79adf64e80cebaefcb119f91a;
// music[6265] = 256'h730de008b20cb21c682b442b5a26f41f31162c0aaa01bb036d0abf18d51b73f9;
// music[6266] = 256'hacde19e902fb41fc48f167f7420a8418981cf90b9101d90577029ff7d6ebaeef;
// music[6267] = 256'habf1fddbacccedd1f2ea8a05a500bdea8ae3aef7f60c7c07a40385090b09fe04;
// music[6268] = 256'h6af9efed1ce558e62afa8c02de0497041fe6a0cb6bd5f7f4fb0901fd13e223ca;
// music[6269] = 256'h31c7e4df8beedeea13e2b8db40de76e2cceaa7e554c745b612b30da5c59c09a7;
// music[6270] = 256'h71b1c3a9c69e6698178deb9aa7bd5ec88bc31cb9d0a911a39fa775b808c1afc2;
// music[6271] = 256'hddc3f6a9c492ac9ad2a943b3c4aa8b99d790309669a748ad7cb675cbafc6feb6;
// music[6272] = 256'h74bd22cfc0d54dcdbfcb85d52cd8c4d294d0c8d86de34ce46fe3ccec78f31eea;
// music[6273] = 256'h04e49bea14efa3f19af440f666f973006e0a600aa9fa52e878e93104cc1b0c1e;
// music[6274] = 256'h9c134815bf28c92b9b21381c291493179d255d364c4437345b16a60e5914d312;
// music[6275] = 256'hfc0a1b16a6385153c95b105d40564142bf20b70922103c14ae0efb1df83a694c;
// music[6276] = 256'h26496b40b33a142c0a231528362d022f8b322640614d15515a57a1613b600848;
// music[6277] = 256'h3434f0367f3b163d913a4634b8346441545d1c6d3f5ef047793ea149615c1b62;
// music[6278] = 256'had54de3ab32b1535184f715eb850693e1d3f7750a365c666f549f42c932f634c;
// music[6279] = 256'hb766cf62814e1b4bdd51385eea66e2574c41ee36d045bd608b695f6c1b73a975;
// music[6280] = 256'h7463bc40e53968445241753c8f3701349434d137873cd636bb29a426d42d412a;
// music[6281] = 256'h2b1daf17e01615164607ebf0f3ed5dedfae5c6e37ae4cce419dfb0dae8daeed5;
// music[6282] = 256'h59cf96c8acc344c6e3cb02cc3ccfdcdd7ae279d5dbc095b13bbe66d3c6d476d1;
// music[6283] = 256'h69d381d2fbcdbdcd1dcf95ce94cf03cea5cbc9caccc98dc8d2c516c8f6cacbc9;
// music[6284] = 256'h8ac79fc461c844ccf9c981c551bd05ba1ebb62b841b208b154b75fb945bdeeb6;
// music[6285] = 256'h449c2f916a905489528985902e96268ec09801c07cccffc6f7c7acc138be40bf;
// music[6286] = 256'h91bfbbc131c499c873c872bf39bb43bf62bce9b60ababbbd9ebfa7c093c43fc1;
// music[6287] = 256'h98aaefa152ab24a78b9db89b3ea7efb69caf18987a8a0b90a49ea5a718adc7b3;
// music[6288] = 256'hc2b50eb097a5aa9c16a751c10ac9f2c091c04fc6d8cc0ed008d08bcc17c653c8;
// music[6289] = 256'hfdd365dfb4e3e3e4dae987ed19ec83e301deb2e4b4e895e66ae6e1ec4af526f5;
// music[6290] = 256'h3cf602f2e9dd08d265d708e083e184e0bfec42fde9fe17f2e6e395e17ae600e9;
// music[6291] = 256'ha4f5c40bca120b109918e426a6322a3a6436f72dc531063bf33fb340e9381c35;
// music[6292] = 256'h403ad33baf3c763f8347cc4df445063dde3d7546de4077213e10f51ad92a8038;
// music[6293] = 256'h5834d11fc918091f621f671abb217e39b245543b782a9f22db342b4bed4a0d48;
// music[6294] = 256'he84a314a1f47964af54f4b4b484c605af863c45c28532a5a7e62a2632e5fe35a;
// music[6295] = 256'h4f5ddc5b2e605c5a923da135414148475743113e3e411d424c4c2462a76c2764;
// music[6296] = 256'hf84c9d400c416c3f303b8e387b3cfa3e814d4966616b2067e561e05ffe5e8459;
// music[6297] = 256'he1662a753f6fe06bfc6abd6b666e5e68a16407655c60f660765e6546c62eec33;
// music[6298] = 256'h754ead5e3b5af456df55bc48042f7c15d50d3d0c7b080a184f2f7833ea2d482f;
// music[6299] = 256'hc7326d259a0ac70371179a2765281b2c0d32452b26264526891ef115ea14341e;
// music[6300] = 256'h8c21da1a6819df150819161699f9fbeec7f867fb5dfe830723194121cf15ae00;
// music[6301] = 256'h5def6efdd11b8423ca11c9f887f1a4fd330ed414bd0602f375e8cde74feeaaf7;
// music[6302] = 256'hd0075f11d20a1b07cf07b8094b0c68071f07af073bfff303ea12d615cb0a4ef8;
// music[6303] = 256'h94efebf6b402c80a1e004de647defbe26edfbadd86d9a2d27bd6b3d9fcd84fd5;
// music[6304] = 256'h01d186d47bce85be2eb42faddabbd1db48e18dcaf4b2feac87bee0cfa9d82be1;
// music[6305] = 256'h42ded5d610d44ed2c9d32fd5c8dc90d84bb962a807abcda8eda682a537a5cea5;
// music[6306] = 256'hb7aa6fb614b9edbbd2c549c5dabf81bacbb92bbf43bcb5ba38bb85b879b681a0;
// music[6307] = 256'h5d8be890d599ca9c5996b88e108a2d8815a19eb9ceb7ecb06daad2a942adfbb0;
// music[6308] = 256'h02af9a9b028a4a8ac49b91a7c2a3f2b467c8c5babca678a0a3adc7c19fc4d0c2;
// music[6309] = 256'h6dc5bdc318c207c01cbf25c229c2afc181b2fc929a8b20a494c1e2c35ca8559d;
// music[6310] = 256'h6ca23399548a5284609340aa92ad67a80eaccbaa9195a7872c919792818b3095;
// music[6311] = 256'hc3afc6c211b7e29fcd94db96fb9c8799d0a34fbfddc64dc200c69fcc6ccd0ccd;
// music[6312] = 256'heacf57bf0ca61fa5d9ac10ab79addfc3aedcced78abf30b580bb80bc80b65cbd;
// music[6313] = 256'head556eb78e589cbbdb96dc378de38ec31e268ccdfc0dbc4a3c34bbe3ec8e5e3;
// music[6314] = 256'h59f56fe667d0c8d5bff2f907410b4a090e075304f2f633e67ae69df7f40b670c;
// music[6315] = 256'haaf9e6e85ae451e769e1c8e6ce038519bf14daf017d29dd6bedc7fd8d5da3de3;
// music[6316] = 256'hade73ee681e5e4e382ea2f013e13a20da9f68ee74ce883e81ae94df346fda4ff;
// music[6317] = 256'h410453105818130f30fdbaf74bfa6ff88afb65046e0532055817b52e64275a0c;
// music[6318] = 256'h2803d10cb91512145b1acf31703b3736cb37793bbc3b6e3bf53d9e361521dd18;
// music[6319] = 256'h8b2099232522052c5e43a35301521d4901457c38151e7118b6247b2668337754;
// music[6320] = 256'h3f662260c85ecd6c0570d155543e9c413f46e141a6436358f46d2f66db545345;
// music[6321] = 256'h063f7d5448661d6b436c1b5acc3fd9295c21fb2e114612507a42122fac284d36;
// music[6322] = 256'h9f4c16514b41cf2ab326a93f2b5bba633856ae3e50349b404852fb53b0476d39;
// music[6323] = 256'h11383248c35ad15949406a2ef22f7d2fc12ecd31d6316b31553d6e53605cf951;
// music[6324] = 256'h223f9233cc32ef30bd317536bd39483af0356b360f3a6b394d397c3a3d3d273c;
// music[6325] = 256'h9134ac2c7228d82e3d38c7385b34b12b6b20ff23f63d12508250734f6440df39;
// music[6326] = 256'h9f555a68ea62d25f1d655e5eb442442f752d3c321d39303fc44d3b5674520255;
// music[6327] = 256'hdb4c0936f828ed262c2aa92f3631c5324235f12c4a22171d95172c1bcc1cda13;
// music[6328] = 256'h45104d14311e1d22c91c4c16840abb05ae03fbf3c6e43deb63060514bf05b2ee;
// music[6329] = 256'h0cdbd3db67f26d05abff93e8a1d954e138fa590462f912f8adff2a04750226fb;
// music[6330] = 256'h66f9f9f8d8f079ef34fab2fda0f958f697ef4fea6ae974ee3ef4e9f473ef7edf;
// music[6331] = 256'h91dd66e448d7ddc877be6cbe7fcd01d211d466ddd2e186df45dafad4ffcf4ccc;
// music[6332] = 256'h1fcca5cf9cd08fd888ec5ced6ae1b3e3a8e9b0e759e774ed63e305ce6dc9cfcb;
// music[6333] = 256'hf1cc9ecbe9c75bcad3ce6fce16cd43c901beadbd7ac418b3079c909ca9b39ac6;
// music[6334] = 256'hb3c2eabc3cbda1bd89bbdeb75dbcc7bf58c009bfb0b6d8af51a6f296b990229e;
// music[6335] = 256'hfdae5aacd4a93cb69dba57b51ab5bab1acaa64aa79b0c0b7a8b4adaa69a4aea4;
// music[6336] = 256'h53ade0ad81af97b480a0ee8870846e8a518dad8a9f99d5ab76ad5cad65af83ac;
// music[6337] = 256'h73a90aba29cc61d001d65dc883ad27a272a2baa756a9b8b7a5d0ecd227cebfce;
// music[6338] = 256'h67caffcdced5eed5f8d007cc4ad29fd25ec14dbd04c1c1c3e3c6b6b19f9c03a4;
// music[6339] = 256'h12b7fdc44bbc11aac39f61a2cbba9ccf00d1b3cd23caabc613c599ca2bc9f5b4;
// music[6340] = 256'h26a909b5dccb0ad8b6ca51b7bdb339c394d86cdca8d813dad2d60dd5d5d787dd;
// music[6341] = 256'hace4dce820edb2e9a9e76fe9f6d63dc764c773c3efc275c6e8cbf3ce11cb19d0;
// music[6342] = 256'hd6d2c3d592eb45f710f2abf020f27ce8d6cc96c50ad73cdc48e6c3f1bce9fbe5;
// music[6343] = 256'h25f061f9fcf858003a1083171c208d26ec24171f471529141c1a10202e1e4014;
// music[6344] = 256'h950be0109a2bba305b1b4f163715af13e417761dd51c57060cf1d3f785138f23;
// music[6345] = 256'h0e16c402c5fbb90c5f28bd321a2b8b203225e729ad25f022781c05160814e21f;
// music[6346] = 256'hdc2b8a24a123182e2f376538ec369c31cf19020cd2123b164d17891f06354b45;
// music[6347] = 256'hd0464f4297412741932e5b206a21ef245a2e172f942da72af9223322b51f0a2d;
// music[6348] = 256'h194c8558694fcb41223de5369126b925453d0e4a0946d551ee60be610863a964;
// music[6349] = 256'he760fb50023fa440ab555e6942620649ec368234c945c8587658664a2e35d823;
// music[6350] = 256'h222942363c3ce544f74797405e3a653c9f3be225ed13d61e8e36883f672d9118;
// music[6351] = 256'hce1a61325145ba400a334623301ce02bf941ff4281276712121434155016d41d;
// music[6352] = 256'h39217e1a3d13bd1428183e17b71207114216421a9d16471b4430c239f931f332;
// music[6353] = 256'h943e193ba9231419541aa8134a128e144914321792151e11a711d711620d8009;
// music[6354] = 256'h710fe2189713bc1481257f2a3f37884afd49884a144b51495a483a409b3fd743;
// music[6355] = 256'hd847ec47a83f2542eb3fe52a6c1bcb1d08318e429533e5126d082f11d11be823;
// music[6356] = 256'h2d294a2f442a7f23da25cc26ff2a462a8c25f723911e701f2a23092ac32c5018;
// music[6357] = 256'h9e006cfbfc0a5f1a2b1fdf26c9279d25d323241cc2186e19e220641de402fdf2;
// music[6358] = 256'h7af26ff4b4fa8ffd90fa90f6a9f8e9fbc6f31df6430a2812a3127212cb0d7511;
// music[6359] = 256'hd813d311bc118f12aa150c0e140ae50c35fb5de796e3e4e445e2efdf1bf29410;
// music[6360] = 256'h6b1d69189b18171e2820d1202c126ef13fda8ae523086d1b9719c01190076efe;
// music[6361] = 256'h4501f90cfb0668ee13e18be9a8ef2ae87ae6f0e24cdf84e274e0c2e4b7e85eea;
// music[6362] = 256'hc4e902d1babc42bee1ce4ce537e409d32fc2b4c1ded7e9e4bae3cfe2dbe63fe2;
// music[6363] = 256'h0fca08b81ab551b454b5bcc22bdb4de677dfd4da33dc5bd4aac50dbb3cb041a9;
// music[6364] = 256'h96aa87bdbcd6b4dc2dde86dd6dd907dcafde30e16bcce2afd8aef7ae91ae75b3;
// music[6365] = 256'hedb2a1b2ddaf03afc8ac83b13cc868d77cce4db8edba2edd08f569f9eaecaad5;
// music[6366] = 256'h5ccca2d85def02f82ee6facb84c54dd79fe761e734db53cc99c723d368e09de1;
// music[6367] = 256'h24e3f8e02ad0dcbde1ac1da959bb5fc9e7c92bc7cbc61cc713c409c4cdbd60aa;
// music[6368] = 256'h699d57981e95799b5ca574a5b09c00977997c3993f9b199898947a94d998bca0;
// music[6369] = 256'h09a402a560a19f98d895dd94ff94d6939a9373a78bbeebba4aa20a8f698f1092;
// music[6370] = 256'h728ef79238a473b53db9f2b4e2b307af7f997e84fb8ceba513b187aeb3b008b1;
// music[6371] = 256'h45a500a3eea8e6a43d9dbe9b4ead02c232bf89b506b1b9b2e0bc95c359c621c3;
// music[6372] = 256'hc0bad3b499a6c69cb0a5b4a9a49f429687a4cec37dca08b96da3bf8d928fdba8;
// music[6373] = 256'hddad3297388b6991a494c98d3d8c639ff2b02fb5b6b832b34eaf1cb61cbafbbd;
// music[6374] = 256'he0c084c086c023c016bfa0bebac506ce8dcd6ecc5dcb08bcb8a5e7a5a3bb4ad3;
// music[6375] = 256'h88dad4c22aab52ab65b1b2b6f5b7ffb63ab918bcdcc1bec257c39fd57de832e5;
// music[6376] = 256'h71d0d5be87c44ad6abdd1ae137ea2ff017ed5ce6bde1e9e57df0a4f153eb29ea;
// music[6377] = 256'h3bec73f0fafffe0b23f9d8e208e16ae3ccecfff3eef362f1d3ed8d02bd173f18;
// music[6378] = 256'hcc17bb10460eb015ce221f24de04eff67ef6d5e5b1e30ee756e451dee6e4f905;
// music[6379] = 256'hfa12e70cff0e1a0ee8100f167917281a4f1dd21bd212e012b717d60a93fa79fd;
// music[6380] = 256'h000fda1eb222c120a127242a0316c4023407c31948272d2a622ede34fa323423;
// music[6381] = 256'h9212e5171f28cc2c8f2dd234043b3e338d2090186a289c3d323fd335f0342e3e;
// music[6382] = 256'h95492f4db149c642f13e6343dc397525f522b423111f0922b03075500762df4f;
// music[6383] = 256'h36405b405d407a3e4f411355046bc7648349a638823f5749cf45de47c45a366c;
// music[6384] = 256'h1f674e4f15426c45793d562d6737a150cf55b450ed513f54d4532e537653c946;
// music[6385] = 256'he931582fa93fd454f359e74671359e36223e0f3834337049055ee9526b3e123b;
// music[6386] = 256'hf24213455940d23cbb458959e05f66508e41a13f713b03332f3f1d5d756ac15c;
// music[6387] = 256'h4e438534a33fae566768146eb96db46fc15b743d713eae4a954efe4de3459d3a;
// music[6388] = 256'h01385b4c9f6439687f5a1e46084253407e3473426e63ef750073455d39497f45;
// music[6389] = 256'h4649d252e961886bc26ec062a14a13445648f14869496b480d471a41804d3b67;
// music[6390] = 256'h685b243e4b2f812ddb3caf48d848b0453241e93eaf334328b52cff32362d5d26;
// music[6391] = 256'ha235954af344d22da21d6f21b02745201720d832db467a3fd525031d79218a22;
// music[6392] = 256'h741e2124a6362a3ef03d524030410232e514c30e5511a80677085812fa15d414;
// music[6393] = 256'h101a1827b928a81c060ab5024d105d2212264711be0112073807d6fff5ff0b0f;
// music[6394] = 256'h971ad417d10d3fff17037e0dff05ad0c162b483f7931e6114c002508a521e930;
// music[6395] = 256'h4a280914d206f40e6f1f9429c12a692b242ba415c3fb90ed18e3b5e400e5c6df;
// music[6396] = 256'he5e01bde3cddabdf5ee4d6f592fe49f1b3dedad311d60edab6d94be056ee18f5;
// music[6397] = 256'h2ae862d3a8cb7ecfded520dc48dce6d5edd0c1cfe0d062cfeacca7ce4ecf73db;
// music[6398] = 256'hdcee47ebedd8a5c64ec43edb8ee779e2d3de79ddf6dc87da45e2e0e85dd44dbe;
// music[6399] = 256'h09baceb5d5ae22b48fc602d6f5d2c7c339bb13b940b518aa85aafdc642d569d4;
// music[6400] = 256'h55e2efe55ddd41dcf7e524ee95eab6e4c9ce28b63db6bdba69beb2c07ebe78b8;
// music[6401] = 256'h6eb431c9cde023e105db32dad7d46cb53c981b9d4fae5cbdacb7359e1a941d98;
// music[6402] = 256'hf59a30994c9b81aaa7b1a4a8529ed795299af2aa21b409b5f3b41eb443b563ba;
// music[6403] = 256'h8eb987a89c94658d8b9d42bb77c3f1bdc1bd93b0f9958184a18d25abf5c3b4bd;
// music[6404] = 256'h29994b84738b4d94f19b779c6794018fd89353a8a6b961b09597af8a8a8d0b92;
// music[6405] = 256'h19933391138d1d8a529353a777af66adedb47abc8baa00936b9b4daa29a6c0a5;
// music[6406] = 256'h56b626d285dcd4c654b049a67ea158a287a522aa10aac9acb4bf3dcb75c65bc5;
// music[6407] = 256'hcec8d8c238a785907d98aea0649db0a269afbab7a4baa5be49bed8b1329e2a97;
// music[6408] = 256'hb8a782bb6abf10aec997fa96f4a610bc2ec4eeb432a8a9abbfae70a5bfa716c5;
// music[6409] = 256'h2fdbb2dc60d8a5d54bd1a9bf91b0c1b797cc38df8adfe0d034c566c663d43de2;
// music[6410] = 256'haee1facdd2b97abd10d22ee50de2fecae3c174c380c0e0c1bec38dc331c4d8c8;
// music[6411] = 256'hc1cec9cf99d12cc933be1ecc98e5dafb9dfe92ea2fe437f184018f0637f879f1;
// music[6412] = 256'h65f707f5a0ef4defc1ef0ceec3edbef2def6a2f647f8f0f7cbf5c4f612ead0d9;
// music[6413] = 256'h1fd906d8aee70105ab06f2ffe8feb9fc1e041f0af80cfa0db30c4e0e3eff87ed;
// music[6414] = 256'hf1ef3df211f2e5f569f76af12eea6bee5cee2deeef048c15a210ad0e1010e411;
// music[6415] = 256'h70163f188717ee10880ab10ff017a51c291d2e1e202118170b02c5f90d0a8a1c;
// music[6416] = 256'h1c19b211c217de211d25ae247520760cebf94902d31a812926241a1de31cf41e;
// music[6417] = 256'h17257429712a0b25e41a8023243d8e48b0451645c6418a42aa48884a454cd545;
// music[6418] = 256'h6340c7449b48464eb5448f3046282627e729fe20481abf2a0d34cc3106375c39;
// music[6419] = 256'h5a2a5717b5135c16db1490179129da3a6f39bf36823e1b426f346c215f182a13;
// music[6420] = 256'hfa11721bce2ef03a313cde40ce418b3fc73ff83ff941b3410344bf3c8828f920;
// music[6421] = 256'he42bf741524dbf3fa627e31aea2c7e489d4f77408e292922cb2f47443b4a0339;
// music[6422] = 256'hd422ad1f07342f470a477435f8230122312fe241e043fe383d2c2427b1411258;
// music[6423] = 256'h7a56dd5bc761a45f985b375e845b2e47ba3bd33a983b4140854192416240883f;
// music[6424] = 256'h7a3f6c3abe3117327e3ac1309a1fcd1dca1e431efe1ba51aa51e161ff31a5e1b;
// music[6425] = 256'h3d210826ab261823e71e3f1c7e1efd24de1f0d20ad301237f037b03ed8443e3e;
// music[6426] = 256'h7e24f013031d2a2fc737803a7d428a44c53a852c5625e42d6538fb39ea35e330;
// music[6427] = 256'h242daf309839fd394b322a2c8d2f5e36df305727f1210520e623ef29632f5134;
// music[6428] = 256'hb5378a3696291f129b05390e2820cf2fb8263518a424912bf2202917221eec3b;
// music[6429] = 256'h4d4b124a764c60472540bf3de63fa0445e44b043b245d04574412c3b9039e83f;
// music[6430] = 256'h963e5e2d2728342f9e2c6528db232d1c901acc233131682c1e16860a590c290c;
// music[6431] = 256'h6c0aa00ca50f76103d19fe2cca33af22a70b6d04c316a62a892b222a7a2e7230;
// music[6432] = 256'hb230952ffe2aef27b4285f284b26fd228722d326332a95293a22811a5a19681b;
// music[6433] = 256'h26215123b420c621b31b950700f8d1fdff0c4916211f2d27fb260f1478f550eb;
// music[6434] = 256'h6cf3c4fb48045302eef393f050099a27f62f342dab29e529522e9a29ff219722;
// music[6435] = 256'h23291630222f7e281e221f1f3f1ff31fa520b42064240d27c51c05094df375dd;
// music[6436] = 256'hb1cfd4d1b2d665dde3f0e5fa75efb5dbe2cdd3d533e717ef20f2a0f874fdd9ed;
// music[6437] = 256'h71cf47c36bd69bef46f451eef5ee33f5e5f934f77df0eeeb0febaeeeb6f49ff7;
// music[6438] = 256'he1f57cee14e5cce246e75bf0e9f06bdd5ecf86d464e2dbec31e15dca62c219c4;
// music[6439] = 256'hc7c2e1c393cb84cb70c4f1ca47de49e45cd38ac134bceebef7bf2cbefbcb86dd;
// music[6440] = 256'h44e30bf1defaa4f4e9f4edf89bfa4ffce5fb43021507c20319fdf2ed7ae8c3e7;
// music[6441] = 256'h76d9e8d698dce6da08d879d349d555d09dc5c7d032dfcbe0dce273e234d491bf;
// music[6442] = 256'h5eb9d7bb9ab805ba0ccb64de5ddbbdc7d5b848ba58d15de6cde76ee3b9df8fde;
// music[6443] = 256'h92dd2dda67dcf2e159e5ede38edfefe3f3e345cf09bf55c98ede21e700e581e9;
// music[6444] = 256'h7df123eb18d7e2c9f3ce68ddd4e53adbfdc5a2c2c9d537e9e1ecc8db73c618c0;
// music[6445] = 256'h9fbebcbd01c41bcc62cf85cf7fdd9fecc3e5a4e071e234e100eab2f822008f01;
// music[6446] = 256'ha806e50285ed9de4f2ebceec1fe64fe954fede0e810613eec9e139e4cde32ae9;
// music[6447] = 256'h73ef07f24ef3a3e164ceeacfd1d56ed043c763d1b4e458ea5bec32f596f736e2;
// music[6448] = 256'h05c4d5c259e007f63cf326e81bdf59e0b5e75fec8eea78d595c186c934e499fd;
// music[6449] = 256'h13f92ede3bcb30c654ce05d5fddc3bed89ed6de619e983eb90eed2f2a0f698f5;
// music[6450] = 256'h96ef1fefdfe50fd27bcb44d402e291e1c2d40dd47dd9e4d599c66bbecacd59df;
// music[6451] = 256'h76e7c2eba5efc3e81fcc8fbb07bf2fc395d6bee994e9c3e677ec3000c20c27ff;
// music[6452] = 256'h99eb80e0f2e8d803dd144f19711ca518f60c0f05fe0aae074ef2d0ec88eb3dd9;
// music[6453] = 256'h16d0c9d31cd4e6d5c8e63dfcb0fb59e879d6b6d517e740f3f3ed75dc5ccb0cd1;
// music[6454] = 256'h6febdafe20fed4f4a2f253ec97d981cfd5cf6bd299db13e51fe588d9a5d975ef;
// music[6455] = 256'hd0fc82ff4302d5fcbfed51ddbbdd81ef83fe48fdc8f613fd5bfd93e96ddb89dc;
// music[6456] = 256'h41da8fd2a3d03dcef7cd61ce2dc9f0c93fcc95cf5fd104ce76da22e541dcd3ca;
// music[6457] = 256'h2fc1fad327eb6ffa0e085d039ffc72f66de851e481e72df17ff9adeb62d722d1;
// music[6458] = 256'h6dd496d8d6d882e2c1f99c0048f1c5db03d315e760ec50d858db0ae869ead3e8;
// music[6459] = 256'h94dfe8d640d4a5db54de75c99fb93cbec4c106c2a3c41bc48dc1b5c65bd71be4;
// music[6460] = 256'h03dc9ccd9fcaf9cd9cd067d18dd2f9d09bcc8ed447e95bf12de293d406d456d4;
// music[6461] = 256'hb6d5b5d84edb63db2bdb8ce967fa56fa1ef61ef637f42df222f5ebf30fe4b7d4;
// music[6462] = 256'h62da63f1a302de01e8fe5c00b6f2d9d767cbdfd20fd956d96de6b6f628f787fe;
// music[6463] = 256'hfa14d91f0214bcfd91f6550037049d06b7131d1e951bbc17f91be31b300c9dfe;
// music[6464] = 256'hc4088420c52bda227d1beb1c7f0ce1f2faedf4f204f3f6ee9df24e07d815710e;
// music[6465] = 256'h62fdc8f1d5f9a90e4a195e0f09fbb1f273fdef10661b3d1095fdc0f99109761b;
// music[6466] = 256'ha01a7a0a58fc8801251763287229b919700a3a08350cf80f531306229e306a28;
// music[6467] = 256'h2217660f00186f25fd236e156b069c04380816056705460ac50e8a0f280bfc09;
// music[6468] = 256'h410ef20d0407790358056f0e04182f14fc0d1109a30d7721dc26fc23d028482a;
// music[6469] = 256'hf52c5f2a45290f3baa4ab446d0377031ef34ca2ed426e126ba26e5276e2bd531;
// music[6470] = 256'he534d32e4c2c432d5b2e3033e036263a92384a30202d8632a73d2544d23e4834;
// music[6471] = 256'h632b232b6d34143af9367f347e34f9363c398c353f389339892b061f141d4e20;
// music[6472] = 256'hec1fd1265b3e67477e407b405c44f9440044b245df3d9f278219af24bc3ea849;
// music[6473] = 256'hf046b148a349ce453f3f3c38fb35203a3d3e103d7c3dfa3f6e3e963f7f47d445;
// music[6474] = 256'h6244cb5037539053384e2332672cae43cd5b6b6da1692f54d9409545605cc26a;
// music[6475] = 256'hc46d8c6a7a671f5a2a43613a863e88446243b149505a945e705fce59104f7c4e;
// music[6476] = 256'h57476b40d9444a4a054e534d8445ae3c073fc84b7b565c56784e76448b300925;
// music[6477] = 256'h1a2c382f9b302232742fc22d7a2c3b2c3d293131f9481551094490350030a738;
// music[6478] = 256'hdf47c44bf83d442d532a093aa94d844ed346cc453b465c4ab5495f44d1465945;
// music[6479] = 256'hd540053f6a40e745a03b2c2f722eba233c13d50e8c1cd529202b282e622fc32f;
// music[6480] = 256'ha82c0f302f3e49344029a2307e2b34229e1bc31a10245429352bae27a71e1f18;
// music[6481] = 256'hc1143025c04133486a458e424b367139733dec2e4726a71e951714184b1c9f22;
// music[6482] = 256'hb817790600035c0055f998f7df06af1bef22bf22d21fcd11b1fb91f170ff1a17;
// music[6483] = 256'hfd1f301f2421fd1ac1144e194f21b7222b1c6019311077fd28f95e0948193616;
// music[6484] = 256'hf814211d361c2014c10d090fbd0fc611bc13e201ccee26ebe4f45b01d1feb1f2;
// music[6485] = 256'h6ee91aed7af8a5fe15fc9df026e9dae214da0ad155d8b9f347fde8026414da1b;
// music[6486] = 256'h9e1f931ef51e41128af58feca2f0a2f26ef1edfd2d170a1bda178f14720da20a;
// music[6487] = 256'he10c9711df04fff3e6e51fd121ce39d44bd782d756d246d132d166d488d79cd4;
// music[6488] = 256'h13d9e4e76cf4dbeda3d430c2eacf2bede9f941f6d4eaf2e287dabbcc90cbcdd9;
// music[6489] = 256'he9ed4bf299e0f6cd8dc9bfdb86ef92f485f6d8f879f5f9e24dcce3c8abdb06ec;
// music[6490] = 256'hc0eaefe70ee6b6e63be825e510e447e074e2e5dff3c8adbd80c02abf50b9f5b5;
// music[6491] = 256'h2cb87ebaf8c449d624dee6d359c1f3b8dcb907c567cd3dcd49d228d20ad16dd1;
// music[6492] = 256'h9fcd74db84f00bf3d6e41bd3a9cf48d6a8d144ceabdc2ee96be978ea35f136ed;
// music[6493] = 256'h78d8ecd10bd4b1c255b024b2bbc372d2ead20bd1d4d100cb7cbd3db811b9ceb3;
// music[6494] = 256'hcbaaa8b461cf35d5c8cd6ecf3fd2c2d534d6e2d452c825b2a9aff0b76bb8b9b7;
// music[6495] = 256'h0ac34ed36bd1ddc115b074b3c6cb58d60adcf4e440ebb6e959d44ec5dac66bc5;
// music[6496] = 256'h8abf16c0b7d306e36ad7b0c206b381b57aca52d957d6aec418b86dc38dd52ade;
// music[6497] = 256'h3edf5ddd75da3ecbf0c150d483e643f1f0f6fbe83ddc0eda8cd391cf07d255d6;
// music[6498] = 256'h58d6bbd781e940f724f0fae0eed33cd856e819f88cfbdbdb39bdefba3ab9d7ba;
// music[6499] = 256'hdac2f1c8c8cb3bca0cc941c54fc744cb0fc754d1b1e745ecd9d9dfc618c162c1;
// music[6500] = 256'hb5c7bdd014d9b2d664cd29dc01f14bf5a5fa5c0347067cf4b8e0c0df37d6c5c7;
// music[6501] = 256'hb1c7dfcd1fcfb5c93dc622c342cfe5e7fbeba3e9a7e866e454e52be02cda91d5;
// music[6502] = 256'h33d485dc4bd43cc0cab888baa1b846b8a1cb76dd73e03ae08cd9e2d238c4ebb9;
// music[6503] = 256'h4bd108ee93f4a1e805d518ca28d50deb31f117f08cf49ff750f855f8bdfb1cf2;
// music[6504] = 256'h78d8abcacad5cfecd2f6affbfffed9eb9ed793d46ddac9da6bcb8ec1b5cdd2e2;
// music[6505] = 256'hc7ec5ae02cc8f3bcd4c824dbb4df37cdf0bd1dc5efcc14d0ffcec6c9c6c5a2c3;
// music[6506] = 256'h63ca87caebcc58e119edceef4af5fff9aef1efda17d2bad7bdd952d6d1dd9bf4;
// music[6507] = 256'h77ff80fe51ff73fc9beb39d76bd82bddc9da4fdaced210d16bd461d2dbd117d2;
// music[6508] = 256'h3bd8eade5ee1b4f09700b2fe28fd08013a028d035f0081002100fcf4abf93410;
// music[6509] = 256'h4321a422920f10fd0400ba12d9215d1dff0bd4029c0ae8194523dc1c110df507;
// music[6510] = 256'h94153c25e81b150a5708ec08da0ab111d9138610ae0e9e0e8501f7f078f44006;
// music[6511] = 256'ha61262130a14371b4a1b000adff82ff5b0f522fdc1043b03cc00c1fe29ffd101;
// music[6512] = 256'h03029e02750508092e0c490f1e0fa70f6c0d490815086508a51690287a280b2c;
// music[6513] = 256'h8e2f732b57250f23fb261e19dc09040f47129d0f960c71140524f523bd13c805;
// music[6514] = 256'hd90a2a1f422ca22b492b8527692398356445bb425c40463eda3d073cd43b8843;
// music[6515] = 256'hca49104dbe484d424441583adc2d322cdd396343e53f523c7d46f04c962f2210;
// music[6516] = 256'h7b0f661c74325f3ac0259012ea0a1f09220db2112a1406137018da2d8238bc32;
// music[6517] = 256'h46335c3169344d40a540b13f8f3efa37b4388d41594ad04a0e495e448033c425;
// music[6518] = 256'ha627302b1a2695250d34e947894b5e36f6209f18d219cc1d421c611ca51bcf1e;
// music[6519] = 256'h23331241533a41316f30912ded212419b125ff3de241383a0a3b483ec5424041;
// music[6520] = 256'h263c6938c93e4056625dfe572b5cad508c3f8e42cd521c635762a550e5454748;
// music[6521] = 256'h5a48cc40f34079534e632664a0652d684c631246d020c9220f3a9d46f240272b;
// music[6522] = 256'hca216926702805208d1bec2e313c893d23401b38c0301d2f5a2dbb28c525da2a;
// music[6523] = 256'h2920080ea50b7d0a5b0663045709590e170f481e0b2ca3243a14c10536081218;
// music[6524] = 256'h2723811e5f0a8b014b0595023601d401b5010b008c01ea12bd1d7613cf04c0f9;
// music[6525] = 256'h02ffb50e3b105e0a190b450d410d060e5e0db6029aee09e7e2f2dd010716b426;
// music[6526] = 256'ha22767253016ca00f6fd2000a0014203bfff99fb89f6eef60afaf500b614071b;
// music[6527] = 256'hbc0ebb0c56161b18720413e8aeda45dcb7dd25dadbd6bed7ebe79dfdccfe3df5;
// music[6528] = 256'h96f41bf849ec17d99cda2ae202e18be0dde8d7f9b4f92be813dcaedc1dee95fd;
// music[6529] = 256'he9fe31fc81f89ef5d5f466fa5dfca0f010e31ce0c5eb88f78bf64deac4db46df;
// music[6530] = 256'h08f059fc0d001afe87fd3bf647e2a1d55fe07cf449fce4f0bcd9d6d2cde1f1f4;
// music[6531] = 256'h9efc02ec1edb96d76ad557d7e9d8f8dca1db81dd6dfb6710380f3a110c140610;
// music[6532] = 256'h71fb91ec86f265f612f9e4f9d0f6ddf61bf5e2f3c7f579015617ea1ef70f0ffb;
// music[6533] = 256'h60eb12e0d6df01e833e533dea2d8bcd239d7c6dd39e250e1c6dbbceabeffb301;
// music[6534] = 256'h31fbaafa2ffef6f194de0bda3ee489f630fba3ee78e223e696f744fd6ffab0fc;
// music[6535] = 256'h7c01c7040403820546ff00ed6fe6e6e784e653e0e2e84affce03f50033ff45fd;
// music[6536] = 256'hc0014b015f002c01aa02880316f37ede0adbd0e3c4f22cfa7cee51e0aedb82d9;
// music[6537] = 256'h17da89d9bad96cd812d4eae05bef59f7160d5d18a712cd1002142e0f19fbaaef;
// music[6538] = 256'heafa220fba178f0bb3fba9f36bfb880daf170719661764130f05dc021812c005;
// music[6539] = 256'haaf272f25aef7aeeb0ed7eebcde915ebeffed60e5a0c120808049d04d608000e;
// music[6540] = 256'h990e420062f616fd7205d70ba905d6f147eb27f030f2b4f450f1e5eaa4e994ec;
// music[6541] = 256'hf3f089f124fd6b120317b4122b12ed10890702f616f11afcc9075a0d960e5f11;
// music[6542] = 256'h7e0d5cfc13e942e8edfdc70cc20bb309020e3c0fa3fc76ebdce82de722e97be7;
// music[6543] = 256'h0ae964f67e052c18cc20851d511da61d561c6e1ac31ee819b30427ffc20b661e;
// music[6544] = 256'h7025a613540375fc57f3c9eb84f0c3fe6402a3fd2df1d5dd4cd8e8d8fbd402da;
// music[6545] = 256'h7aed28fff9f73ce087d104d8a3ec15fa49fbabfbaafbebf0dbdb92cfe8da16f4;
// music[6546] = 256'hfd0497088609a50734f596daadd333dbcadf4ae3a3e452e158de2aecf1043d07;
// music[6547] = 256'h10f524e534dee8db76d990de9ced57fd6bfe0cee6be399e15bdc89d717d95adf;
// music[6548] = 256'h91e1f6e3efee84f6c8ef15e09fd7a8d8bed637d6cce09df46308070b88f632e7;
// music[6549] = 256'h19f7810eec122c0d3f0a870ac3fe51ef77f460fb27f567f161fd62129c126500;
// music[6550] = 256'hc9f21ff1b7f8f8ee96dfc5e811f3faf5e3fc9101e9f7e7dd55d00dd7afda89da;
// music[6551] = 256'h6ae161ee77f4baebf0e0c6e01ae3badbedd2bad503e087e544ed03fe59024af1;
// music[6552] = 256'h46dee7ddd2f03f014c00a2eee1de49de8cdf25dd86e228f75d0662fbdee98de1;
// music[6553] = 256'h08e61bf5e1fca9f408e3c7dbb4e4c4f3a001a8fc75ebafe1ebded7e039e128e9;
// music[6554] = 256'h77faf3ff7afe2402150316f499dc65d80be698f07df4b6f724f888f48ff326f0;
// music[6555] = 256'h9ef0bb029516ad1991082df8c3f7cbf486f0c9f149f59afa2bf69ef1b3ee0fe1;
// music[6556] = 256'h74d9c8d5ccd2a4d966de8ee690f640fc67f1e1deffd5c3e00bf6eeff2bf5e1e2;
// music[6557] = 256'hccd9a9e557f683f967f9bffbd9fdb9fba6fb0ffe74f0a8e28ce205e0aad9f4dc;
// music[6558] = 256'h72f3ed0269fc8af80ef8bff8c1fab9fb8e016b024f003ffe55fb2400c2f574dc;
// music[6559] = 256'h78d62edbc6dcf1dfefdedada6bd753d6c4da63dc3edddcdbe0d628e8c0fe8ffe;
// music[6560] = 256'he4fd4901a7feaff4adeb71ee2bfb761363202912f40262047f164b20b81cfc1f;
// music[6561] = 256'h8f25882a5b281721aa1e9b1d3424851d0d05d5fa2afc9001bc08990a3f0a4b0a;
// music[6562] = 256'h400887ff42fdab045e0af50d660151eab6e728fad70f9114380117f02aee73ec;
// music[6563] = 256'h58e9d0e642e88aecd5e9ffeb62ed91ee4c02440f88104813a110e90af3021206;
// music[6564] = 256'hb008a8fe37fce2f9f4f3d2ee23f51010fc1f0e1f8417fa0edf0d6b122f1a5010;
// music[6565] = 256'h74ffc2fd55fb40fe7e03d30144fc08f979074d145d13ff14581f6d26d21a4819;
// music[6566] = 256'h0c1fc00c82006d081c16e420711f061ecc1e63136b0160fbee08cd1de724a915;
// music[6567] = 256'h50fde0f23803c818c01c2a140c065dff5cf99ae4b4dbe9ea80febd065203c200;
// music[6568] = 256'h68fac0e93ade0be673f79efbd2f371f1abfaf0fe60ef1ddf7dda91da44e2aaee;
// music[6569] = 256'h10fb8f02c9f8e8e739e344e3f8e01ae035df24dfbdde33de77df28e2ddf1bb09;
// music[6570] = 256'h0a103bff16e732dd0ee0fedd98e035f42a089a057ceff7de1ddf60e41ee4d2e9;
// music[6571] = 256'h41fea00a4b00a1eb88de4ce5e4f8bc065aff63eb29e9e3f7d0fcf6f78d017016;
// music[6572] = 256'h021d84192619431c402162230924261abc0672ffd2ff41fc71fae10703215329;
// music[6573] = 256'h8b1d8f08a5f49bed3fe824ebee01f113ce0e74f9d0ed12f356f444f121ef00f0;
// music[6574] = 256'hdff635fb3ffb59f524f57a08b314a40c3efe73f6da028c122e16b1161f183b1c;
// music[6575] = 256'he1140affd8f6d405171c9723fe1357fe67f6c9f705f663f9660b87201c233812;
// music[6576] = 256'h680229fc61fe06fe6f006a13251df7174c18cc1d82226c21fb1fee15f0014dfb;
// music[6577] = 256'h41fece027e06a209b80998ff830866253f32322da01fe916131554129f13ff16;
// music[6578] = 256'he816b91709249b35f5375c29d519ac17b31896134b15a12a4341b132590e18fb;
// music[6579] = 256'h47fe6e13d41fe01b931d4722ad1d590c8bfe5804c312241c2e1c431ce2205c1d;
// music[6580] = 256'h240f1804dd01b6fd4cfbac070e187a1e192033259c25e11626059f014a041500;
// music[6581] = 256'h80016114a3290b29781193fd87fbe4001f032c022e02e203130d391f502bec24;
// music[6582] = 256'h5b10d905d211701bad162514c41ca52d8130711fd6187d22aa313438f929941c;
// music[6583] = 256'h111a1e28e845724b3d3508220920393242463244d02c3b1ce31f322663236122;
// music[6584] = 256'h6e315941844519475a48fa439a34052c322d4222de1a6c23c132293ec6373327;
// music[6585] = 256'h3120d3245025aa233c272d262528672c732dd7300f3208331532ad305d34f534;
// music[6586] = 256'had35993459302b304f2e9932694711581f520e3dcf2b852e36423c50bd489631;
// music[6587] = 256'h0f2151246c366046a845753a8e30f82e2828e5116b11cb286531032f092cb024;
// music[6588] = 256'haa219926b72a452bcf297927dc28a6289424b01f401c7c182d10841b972fbf20;
// music[6589] = 256'h8b0c050ced0c0211f713dd10a30f1310b610290e9009bf09a90768044e082108;
// music[6590] = 256'h920c6b1d2627ec1f320100e8aaf4c3069e0607009fff8205d707ff05b2fe50f6;
// music[6591] = 256'hd3f3cff703fdbbfbfcfa45fa2ff906f7b2e4ffd267d5e4e4caf18bf262f635fc;
// music[6592] = 256'hdef7b5f172efc5f1eaef82ebb2eb64eb70ef81ebd8d784cf5ed1b7cff8ce7bce;
// music[6593] = 256'hd5ce2ad10ce01bf8c4fbd2f208eb21e0f3dec0e6ebef53f397eba4e220dbe7e0;
// music[6594] = 256'h39ebd6de37cc0ac7ccc8c2c849ce74db66e087e735f14df406fa7cfa35f86bfa;
// music[6595] = 256'h10fc63ff91f6afdf4fd554e14cf2f8f85bf86cfbc9ffc2f51ce1cfd732e579f1;
// music[6596] = 256'h00e343dbc6e4b5e3bfe2cce685e8c4e432e0b4e1f1d3aebfeac347dd45f43ef0;
// music[6597] = 256'h31d70ebf97c01ddbf9e7b6e410e0bfdcaade20dfb5e34be3c3d308ccd4cd76cb;
// music[6598] = 256'h99c853ce61df30eb59e4b4d51bcb69c624c689c77cd44fe7f9ea62ea9fed34ef;
// music[6599] = 256'h26f35ff582ee8fd6a6c111c6d1ceffd185cd0dc268be5cc1bdc80ccacbca85db;
// music[6600] = 256'h8ee36ce115e2bde059e4c1e163dbc7e481f518ffa5f30edea8d6f8dabbdffedf;
// music[6601] = 256'h32e61af39af4a5e8f4d830d6f0e784fcd10098fc87fec1f07cd18cbf3ac0ffd3;
// music[6602] = 256'h94e766e50ae1bae135e1c4df2ddf24dda4ce63c20fca00dc02e9cddf5cca63c4;
// music[6603] = 256'h83c922c83fc145bf91c197c430d144e5c4e8b5d509c635c8a5d4d7ded5dd4edc;
// music[6604] = 256'hc9dd59db6de646fcb7fdbaea63d904d8cbdff1e177e7c2f408fbe5f828f9cb00;
// music[6605] = 256'h04ff6ce963da8bdbd2dcc0dc3ddda3dec1df62e59cf69d00defd35ffb7fcdcf3;
// music[6606] = 256'h58f5f7fd72ff49fa12f72dffc4114c1a73154c14e1122f0780f97df68cf847f6;
// music[6607] = 256'h70fa3e097a17331657043bfbacfe87ffa802070138efd7df1ce599f5bbfd21fc;
// music[6608] = 256'h91003a0a1106ecefd8dd05e6b1fd5f0ad50226f0dfe51aed0ffe16075ffd2fee;
// music[6609] = 256'h26ea59f7c005a4ffcaedb8dd02dc8dead4f6e0f5f3e456d952e00ae543e626e5;
// music[6610] = 256'h21e0ccdf47e1aee154dd93dac8e2a6e951efa0fab1ffbbf54fe7dce3b7e6bce6;
// music[6611] = 256'hfde8bfeb28ebc6eb6beadce56fe4aae3a0e491e868e84becd4f7acfca2ff6804;
// music[6612] = 256'h2102f0fefdfe9603ac063303830e471e0f205320b11ab215ee170f198f1c151b;
// music[6613] = 256'h641c801acdfdcce40de688e8aee204e900ff8c0b520bb8080c05cc037107ec0b;
// music[6614] = 256'hc30bae09a607a9063c065f048d07ce0c020f5f0bc4028000d8022408f10815fc;
// music[6615] = 256'haff0eaf49507a112410d3509310a2c0cbd09d20a9f0bb4fe80f8fafe6b0bda14;
// music[6616] = 256'h440967f7c6f032fe38132217d3146112bf0b070aaa0c8b0fba12ae1429147b16;
// music[6617] = 256'h97179b176d16570de7091d0ad40e8c20bb21d9147b10ae0e4a0add098917f526;
// music[6618] = 256'hbc2d70316e32a02a8c14fe08a70c4d0dd110ca12c412fa0e2f0a800956fad2f7;
// music[6619] = 256'h2a0c7310a91034158a137310f60a9909870d7310a212df12f0136f130410e812;
// music[6620] = 256'h1015ec0555f152ef6201171511173f0705f773f49700080e2b0f65021cf257f3;
// music[6621] = 256'h4b066611ee0f960dd00c120dd210ae17ee12e60159f97bffc20cd111590fe212;
// music[6622] = 256'h1d161619381d4d1cb91826131b0ef10a6011bc1b57117efec1f431edfdecf8f5;
// music[6623] = 256'he9fab0f5edf6d90992186a17d1150714e90e7a0a17053a0c7f1e0428ac2c1c2f;
// music[6624] = 256'h882f86221f09af02c608740a1008f30dac22741f7c0df00ae2078a06230aac0d;
// music[6625] = 256'h360d5609f406e5fc1ff6c8f653017e17261fc41edd20e61eba1dea19cc169416;
// music[6626] = 256'h841bd4229a22c521a51b670964faa5fd4c0f5e1d9419e5063ffdb007451b2f22;
// music[6627] = 256'hb31259034dfeb00a561f27222321d6218c20de206621ef2300169205c6056907;
// music[6628] = 256'ha106a5053112171e4d177714c61312145717471ac41e152013230a1ce10e2e15;
// music[6629] = 256'h421f3921f01fe71ba0176e18cb1b881c521f52236726262694249223a21df828;
// music[6630] = 256'h033fc244e1438e459144962bb30fa713dc1ff72b312b18186c0b3b05010c2b18;
// music[6631] = 256'h131a281ade171d11d80a831026146d03c4f32df50104f30c350c8e0d2809cb03;
// music[6632] = 256'hb904b009c90fcc0d8207e2005effe3026dfba0e98ae20df0c703f30a01fed2ed;
// music[6633] = 256'h0bec7fe987e5eae753ec77ef7bec43ebade98cea23fb2207250644035d048f00;
// music[6634] = 256'hfdedd7e340e585e3dce373ece0000d097afd21fe6f0fe81b5e199d162d15fa10;
// music[6635] = 256'h8714020de8fedffec7fcacfa59fce2fd9efb24f579014312391388118d0d4410;
// music[6636] = 256'h2710e10293fb41ed70db7cdf01ef42fbeaf585e180d67bdcf6ecfdf7aef31ee5;
// music[6637] = 256'hb8d866e008f31ff988f748f639f4daf3a7f459f4d1ebb0daacd413e19ef152f9;
// music[6638] = 256'h54f749f598f27ae610d80fd97eec6dfe4602a201a802abfc14ec67e032dfaedb;
// music[6639] = 256'h1fda59def5ddcedde3e1a5e30be27fdfc8e1cee217df7add5ed9e9df4ef4bdfb;
// music[6640] = 256'h0df839f69df78ded58d823def7f15ff3a5f47800e310f514e00385f285ed10ef;
// music[6641] = 256'h20ef00f3a202d20e2508a7f620eb28f12806b00e240a950bb1ff42ee99ed8def;
// music[6642] = 256'h2bf2c1f261ef47edd3ea9fee99ec11db3fd065dc2bf3a0fabeec55d7a2cc68d7;
// music[6643] = 256'h9aeba4f258e2c2cd06ca70d09ed197d03adbe9eb24efa2de93cd53cc43cf30d1;
// music[6644] = 256'h13d21dd360d5b4d9d9ea43f3dfe8e5e593e8cfee05f2c1ed7eeaf8e571eaeee8;
// music[6645] = 256'h29d9d8d71ed926d53dd4a3d111d2c9cf3bcdfdd072d21cd636d6e3d05fda4ee7;
// music[6646] = 256'h45e996ece7ec92eb06ef41eb80eb9cfb88083b096e06da046dfd06ecb4e179ed;
// music[6647] = 256'hd6029c137b17ab0b39057d0b14146e16260583f010e9deec72fbaa00b6fbddf9;
// music[6648] = 256'he1fada00a403f0004bfa58f518f6acea7ddc5edcc3df6fde96dfeff0f0033501;
// music[6649] = 256'hdceec4e099e433f5ef05270432f3b6ebbaec08ee64eda1f42409d81352167c1d;
// music[6650] = 256'h61219316b7020f00690ac60b7309b113ca27fa2d0d2b562bbe284928052a872c;
// music[6651] = 256'h7c252d11050ae6147a29a234a52275110511df13ca147f0d410fd51d1b239a25;
// music[6652] = 256'hd42673291b3a1942eb3532261921e129d42c06271e1f0b11240b4b13a3205c25;
// music[6653] = 256'h7e16b3058c0017021f07810d430dd609be0a3bfc40e7c8e536e74ce671e423e2;
// music[6654] = 256'hd4e3b8e6aef7cf07d0079b089507cf07e509060bf107cef18ddfebddd4df29e9;
// music[6655] = 256'h9fef1cee7ce833def6d9a7dfb7e8c7ebdee7c0e344e064ddd0dce5dbf0da2be8;
// music[6656] = 256'hbafdaffeececebdbeed9e0ead5fb0ffe94fb64fe2efe69f133df81dc2fefe4fe;
// music[6657] = 256'h47ffa2fa50fd9ffef8ee50e1c1e184ec7d00250ca7115117e816a4135f0e110e;
// music[6658] = 256'h8c129713ca10310c100fef1257121b10e30194f2bdf21ff6f6f148f0adef3ce2;
// music[6659] = 256'hc1dc60ef0802ce027ff11ae0f2de82e13ae015e6d2f51c0101f9dae708e260e5;
// music[6660] = 256'h5de753e6d2eb3bfcad04b5044009c208980381013603f205c1025a010004ae06;
// music[6661] = 256'h150c4a068af4cfee4dfacd09210ea408fa0d3916cc0900f875f1e9ee12ee3ff6;
// music[6662] = 256'h000d8f22791f4e0671f2baf54bfd41fc8b00e50d6915160e42010afb0106f317;
// music[6663] = 256'h8b1ae3176317491d2829c8294e2d063515344733d925ee12dc10cd144014ca13;
// music[6664] = 256'h971df12cb52f4f226d12d711572100300a30c922050d85fb72fa85fa1dfc270b;
// music[6665] = 256'he7180817530622fbcefcf3fde2ff3401a1ffc6fb1f011615771bb0155417a61b;
// music[6666] = 256'h811f2a1dcd17870c8ffaa7f925092b19551d710d70ff9302df072103b4fc83fc;
// music[6667] = 256'h07fc8ffbbefec0fd8dfbd808671d6e1fed0f5e01e6fd6afee3fbd70288152b21;
// music[6668] = 256'hb31e421cce1dea17f70963fe9906f61c10283f27a3200e1f9c1da10cb50a8921;
// music[6669] = 256'h202ff82d5d297d226c201a348848b245d43d7539a7390d3cd03c6c3bfb2cb624;
// music[6670] = 256'he928f826a31ffc198e2bf73d0d29920b95009007661b87292123ce0d8801e601;
// music[6671] = 256'h7603ea02ce0613173d22df1df2104106cb0d591a621def1e97236623a31221ff;
// music[6672] = 256'hfcfd190eba1f6b21141b3d1b9f19830cd4005106a915ab1f0a18920233f9dfff;
// music[6673] = 256'h9305ee07df074202d1fd50ffaa01dd026e079912071af6119d0598036905ab01;
// music[6674] = 256'h23012705f9fd72f086f52c092c0c9cfc21ebede0fdeb86feb30648124c22ba23;
// music[6675] = 256'he0112c010ffcc8f93afa8dfd880021fb11fa890a65158e1590125d1144149f11;
// music[6676] = 256'hff12e20552e52adc16e069dce9dadae306f776fed2f9abfbaaff70f717e73ce0;
// music[6677] = 256'habdd64d857da6dea6efe0bffafec0edb23d69fd9c0d74cd9d5e7e7f23ff1f5ef;
// music[6678] = 256'h08f38bef75e284d739de3bed3cf2d1f0d6f019f593eec6daaad24cdc21ef5df9;
// music[6679] = 256'h45eee5dcead662e313f5defa13f079de92da63e609f7b3fd9eefb0dc8cd51ad7;
// music[6680] = 256'heed7d9dcececa2fdeffabbe570dfdeedb6fc1a0a2409f8f8a3ef18ef70ecf7e8;
// music[6681] = 256'h2ef22a073a12ac06d1f125e819e848e87fea53ef8aeedded48ee12e09bd3aed3;
// music[6682] = 256'h2ed19ed14fd5e8d7a0d875d403cf63cc0dd809edabf232e4c9d5d9d5c9d7f4d6;
// music[6683] = 256'h28d709d717daacdb2bdcc5dad0d969e39fedcceeb8e533db29d85ad45ed3adde;
// music[6684] = 256'he3f1bdf6efefa0f25af068ecb5ed9feb22f3d1f96bfbd3fb0bf691f55af493f4;
// music[6685] = 256'h2df55be65cdbe6dc6de211e155dd79ed43fc2bfd37ffdbff050100fdc0f909f8;
// music[6686] = 256'hc7e3d6dccbf040f673efbdf5360a8918a50d42f8f0ec29f3aa03f409d209a40c;
// music[6687] = 256'hf50a8509410c310da60d610c430a330ea80da5fd69e98cdb1adbc7e896f5d2f6;
// music[6688] = 256'h3fe978d6dcd644ec8dfd3bfd4ef6f8f27aed58e0f6d6dddcdbea38f557eff9dd;
// music[6689] = 256'h13d827d9c3d868db45df02e1b5dafede45f032f4e5f54bf91bf8def8cff6fbf7;
// music[6690] = 256'hd3f4e4efb1f3b9e8c7d9b6da11e459eef4eb94e821e85fe3f7e7d8ed63f6fe0c;
// music[6691] = 256'he21c071315fa29eee5f191f624f728f2b7efd5edabf4550a3d10e20f661ee423;
// music[6692] = 256'hd21c3011680a9016cd25192ab026e7218a21d120ae22fe2408185b03b0fc800a;
// music[6693] = 256'h5a1bc91d761cac1c781090035d08e908b3f98defb0eea6ee35ea39f13a0b7116;
// music[6694] = 256'h62121a115c0ec108b8f81deeb5fa2310441fb11835079afd29fd0f0382086a16;
// music[6695] = 256'he1242c236c1f3f22cb252219fc051005260af8094d0a201811230d13a909960f;
// music[6696] = 256'h8c0c23000df019f0f5019e0d94087bf8f0ed60f25e01b40ba105d8f80ff29af1;
// music[6697] = 256'hf9f294f457f3b1ed72e6e5eadefdce0205fa90f947fded088918a319010ca5fe;
// music[6698] = 256'h3bffc009ea116f0ec90056f8f1fc9309da124b106901c6f8f7fb82fbaefe54fa;
// music[6699] = 256'h45e6d3dfc5e0e8ddbbdee7e464ebf5e7e0e8aaf397f9ebf9f3fa8a0189fb3fea;
// music[6700] = 256'h7ce3e2e1f4e403e9f5e883e805e329e022e5a0eef4f4d2f02ceb2ee66ee5dae8;
// music[6701] = 256'h1fe688e139e0ece41de801e82df5830006ff0cff31fedbfffc0557087e06ac00;
// music[6702] = 256'h69ff40fea8f1a2e854ee2aff9f0b580513f99cf328fa7f06fb07e706f00be50e;
// music[6703] = 256'he20e1b10af0f080dd91770261f22401e9f24ce273b28fd226f1a7919fc19f510;
// music[6704] = 256'hd907550f191f0722451d721c3f1cf41ee3218423a8206904c3e7f3e8faeedef3;
// music[6705] = 256'hbdfa36fbcbfa9ffa07fbf5f72cfb7b0b0510540f5c13f40e710c4c0dab11171d;
// music[6706] = 256'h8d212d20d418880f151091106e131514d80314f8eef910fbabfacf01fa12fd1a;
// music[6707] = 256'h4915ff132416c212eb08d4ffc8045d127a16fa10500fc6157a1be51bdc186f0c;
// music[6708] = 256'h80fd14fea00cdc1b6e229c2487263722f91bc717c317601a521bea1d121c361f;
// music[6709] = 256'hf72db22ab31927173c219c2c0d2e9721c4140612cd1aaf25ad1f41110b0e4b10;
// music[6710] = 256'h98119a0eda13c124a32b332d702ad51a9906ebf2d7ed1df728fe87000a0a9616;
// music[6711] = 256'he512c60e6b14c817fd16f60e380c8a0d5810d212bb018cf7d7fafff82000ee06;
// music[6712] = 256'h480c8c0f93068806ee0ca210dd150b16131d922d9a3102266f13960771118825;
// music[6713] = 256'h182f6725900edd0153095e19901f2f16f2097106261262203624ca26092ba42d;
// music[6714] = 256'h962b792d1533d82a3c1fc922d4314b394b3508356d362b413d507b51bd4f4950;
// music[6715] = 256'h81562857e84604424948e448854638412d3d0d3e7f40f34243456147bb496c46;
// music[6716] = 256'hdd412b472d415230c428bc285a372d45613f0e3532329b35d9306f2bac2e4d2a;
// music[6717] = 256'hf81ecf1ab12a2b3edb3fd23e4a3a3329b61b1e1f6222a31451099d0ce316891d;
// music[6718] = 256'hd11c051ce71aad191f121f09660db80df507e705bb04a4072b07d404f3022bf5;
// music[6719] = 256'hd6e60de83ef6bb05d807a4f94bebeeecc4fc2d0b6e0a9df9fbe75fea60fd3f09;
// music[6720] = 256'hfa06040127008ff82be651db62dd25e9aff14ef9550a7d0af50267044dfeb3fd;
// music[6721] = 256'h9a0088fdcffb75f7bcf8fafa01fde801cff2e0dfc6dedfde6edfd0dd77d141c8;
// music[6722] = 256'h4ac874c904c951c5c2c006c0eabf4dbeddbd86c64ada1fe581d9a8c6a5be23c6;
// music[6723] = 256'h7ed6b6dfbad9b7ca7ebf97c81cda15df6de2a0e415df74d9bed43dd5c6d70ad9;
// music[6724] = 256'hb2d9bdcd6bbee2beadcecfde70e0a7de6edf8fdcf2d97bd677d5f1d84cdd36e1;
// music[6725] = 256'h4ee1f1e45de5eed783d1cad2cdcc00ca27ccafce83d3ffd37ad4fbd542d2b4d1;
// music[6726] = 256'hb0d0a9d4e5e939f99af89ff6e9f9edfc27fca0fbb7ee37db98d86fdd0ee0d9e6;
// music[6727] = 256'h55f64cfe6af792f4e7f4caf81ffee7fb7cfb08f2fde44be370dab3cddfd022e0;
// music[6728] = 256'hece85ce8ebe9b1ea04e9e4e9f5ede2ec0ee807e8a3dfc2cf4bca1dd3bce1a1e6;
// music[6729] = 256'h32e65deb86ef8be719d7dbd0f9d83ce64bec0de4e6d4e5ce25d917e2cae6a9ee;
// music[6730] = 256'h9df33ef5e7efeceb1fe6e2d513d055d437d6d3d322d775e6e8ecf6f04ef737f6;
// music[6731] = 256'h1df770f905fc1af3c1db38d228d6bfd7f9da25e9b9f956fe81ef88dd2be672f4;
// music[6732] = 256'hd7f2caf09fed0ceab3e846ec1cee1bed4bfa1f065005ec041b08bc079af81be9;
// music[6733] = 256'h9be7d5f61c088905c9f533deedd9b4ee8bf5c7f1cfeb72f358042dfd21fc0c0b;
// music[6734] = 256'hf2158a179d043af821ff7e055702d5f7acfe680f631391168e1a4b19d1160016;
// music[6735] = 256'hc116d20d5dfeccfd830ad813640e19fc2df691008f0775073a0345ff8efc61fa;
// music[6736] = 256'h58fbbffc8904d313fb19650cb2fb9dfd5c069209300b800a120b6a0acf0e751e;
// music[6737] = 256'h8122b5161b0917047013422529284425b720e11fac21e91ee21d311d9d177516;
// music[6738] = 256'he61ab41b9e1f4b288b29032b5f318f335530fa2bc12d402b4c1e3f166915b915;
// music[6739] = 256'h2412870bd7039cfabff7b5f8a2f7a4ed91e0bce196e5dde35ce07cde6ce17ce0;
// music[6740] = 256'he0e86ef5cef147e9d9dedddcddead3f6b0fab1f955fc33faa1e852dab2de7ff0;
// music[6741] = 256'hf7fdc9fef3fc9bfda4f69be499dc40e982fe620726fa35e750dc6de2faf3b9fc;
// music[6742] = 256'h00f7f8e30edb84e9f4f70800110310042205d8f995ed17eb7ce79ee58fe7f3e8;
// music[6743] = 256'h34e985ebb4f939052dfc41f5c4fc7e05bc073d015fff5309dc11e40e610128f9;
// music[6744] = 256'hd7fa19fb24fc3bfc71f704f69bf659f7aff98cf964fc6efd03f234e614e5a9f1;
// music[6745] = 256'h5303d1064bfa10e8f1e075ecc1fa3ffff8fe3d039101caf156e59fe4eae757e9;
// music[6746] = 256'hcaed21fbae05d000dbf284eacee9ade855e568edc900bc0506028d05f8064d06;
// music[6747] = 256'hc202aa01e50331007a017706660b7d0d0cfc73e7d9e1a7e468ea29f023f602f3;
// music[6748] = 256'hd8eb57f5fb0396074cfffff098ee44fa5b07730ad0fe72f509f545f2d9ede9f4;
// music[6749] = 256'ha2091d12fe069ff6cde876efdeff2d0e1623ea2afb24891fb41b0421e2262c2a;
// music[6750] = 256'hf6280b16f0ff990059135b2171237a213f246923b6128f045002e7046e01a7f2;
// music[6751] = 256'h7cefb1f224ee24edcfeaa5ef7bff9c06c000e5f4b9ef3af13eee5fe889ea34f1;
// music[6752] = 256'hecefdef400005302a1058508590a160b300b5d10cd03e6edfee9b1eb0eec63ea;
// music[6753] = 256'hccf1e8039907bcfc31ec2deabbfd6d087b0feb0e17f6c2e96cee42ec06ef51f7;
// music[6754] = 256'haffb11f932ec8ce73ef5e201270199f888f426f4abf24ef762fd4902f0007af7;
// music[6755] = 256'h97f777f7a0fa0f0d2111050edb10f40f5312ce0e070c6517431ede1a8f166818;
// music[6756] = 256'ha31b9d1ba21c54198111540a290bb817b61c7c102b01b6ff6f0d90107e056e08;
// music[6757] = 256'h3a14f7161b165916e51aa41d64174c0d9f07af13eb1f421bc41893143b0f8512;
// music[6758] = 256'h3714c911940768012108e30af11155225f25b21647108919171cd81a2e204925;
// music[6759] = 256'h1723ef15f80f8f13c415b220c327be22391d7418c51c682677319f36972d9733;
// music[6760] = 256'hba38aa2d423938450044083fad28aa22942d62324e34d327392eea452541753f;
// music[6761] = 256'haf460b399132093cd8398d2fc42e6531b92ef82bca2c85304530cb2d71398437;
// music[6762] = 256'h1220da25c12a9a160816e20f65029f0b8517d31eb11a49122d0c06057d0d030b;
// music[6763] = 256'hdc015f0a000849025cfb18f2f4f6c3efa7ecb6fc6aff8204070a6ffc05faf604;
// music[6764] = 256'h520525faa7f3adfda305130a2112830f190e7d0da104af00faff64092314580d;
// music[6765] = 256'h8c07540a5a11e118ca1e0e24b51dac18241fd7221c232224de28262cd92b722d;
// music[6766] = 256'h6929ff270d2c8827862eef47bf4bd23cf03d5e43a042a043a64306469e405337;
// music[6767] = 256'h933b5d3e663eba3fd738b935b238cb366236273b43369427d2221726c623511f;
// music[6768] = 256'h981f211ec119b81ca523fe252d1eb8162e1f7c20e81451161b1ee61e8321c71f;
// music[6769] = 256'h3b157e1d77279418c016aa1ddc1e6524c31f7d1cbd14c60898131117b4106111;
// music[6770] = 256'h010dbd148226e4234e115d04c1fc5afa4103940c7617cd1c2210fb07b50cc20d;
// music[6771] = 256'hea088c0b8216f21af01490082300c902f00a370cb4096a187329472c7728a922;
// music[6772] = 256'hed279f2d452daa2b82200e1de4189d140a2586284a237b294224f11c39177a0f;
// music[6773] = 256'h820e7305bc00b10bec043ef2f6eb4ced46f068f3e4fa7bf941f033f30be950dc;
// music[6774] = 256'h66e943f03df16efa92f75af49ffba3f4c2e9fff29ff816f13fe675dfdee08fdc;
// music[6775] = 256'h57dd37e37fe025e3c4de14d61ed3d6cb20cdcecf35cbc7c8bac65ac6d7c339c0;
// music[6776] = 256'h37c01ac47dc36fbcc9c5e2d01dc881c354c74fca9cc885bad5b21bbcdcc274c4;
// music[6777] = 256'h00c22dc266d39cdf82dd5bd7b8cb67cab2cfd5d2dfdde7e67be22fd43ad19ed8;
// music[6778] = 256'h17d815d876db65dff3d73ecf3edd95dde6d564de17d753cdf2ce4bcb05c958cb;
// music[6779] = 256'h8ad390dd1be21ae03ada46d590d032d45adc9edc5cddb0dfffe1dee2ffdef0db;
// music[6780] = 256'hd8d4c7d23adf43e2a4dbf2da78dc91e246e7c0e69ee8a6e1c7d50ed999e541e9;
// music[6781] = 256'h15e3afe84ff3a7ec72e773eaa7e6b1dcb9db6ceb29ea8fdd4be822ebebe6cdee;
// music[6782] = 256'h9bedd4f14ef782f0cef10df4bdfe3d0cbefff7fcf20a8a0dc7155319750efe0a;
// music[6783] = 256'hce064704eb0e3917be185d158b0fe90f2a13c418b2178e009be793e087e4c2ec;
// music[6784] = 256'h4eec09dbf7ca44cff8db6be0d4e236deead538de25e37cdbeade51e38ee16ee7;
// music[6785] = 256'h75e986deefd7ebe088e922e32ee1eeeb97e80dddeedf82e1a8dbd7dcdbe15be1;
// music[6786] = 256'ha8dc65df20e8a7e9e6e956eab0e525e89ceb80e634e457e0b5db2dddfce0f2ea;
// music[6787] = 256'h13e7d8d9c8e1fbe503e501efa8f094f2e5f55ff442f9a3fc3efda9fd34ffca08;
// music[6788] = 256'had0f540d9e087c0262029b0b3909e001fc070f08b30964107c0c7b0825f7b1e1;
// music[6789] = 256'h63e276e8deeda8ec0be792e72ceb8ef054eb77e4b7e514e312e33ce538e913ea;
// music[6790] = 256'h5fe7a2ef12f1e1e671e178e2f8eb58f25decafdfb8dd14ee05f6c8ee49e949e7;
// music[6791] = 256'he3e40bde90db4ee4f7e8b7eb66f2eeeb10e3abe356de76dc38e371e898edc3ec;
// music[6792] = 256'hb2e2c5db9be333ec88ead8ed5df164ecd2e343e1b4e517e67ef66e11aa13990d;
// music[6793] = 256'h690e1a127810c406de048a02c000120bc80baf05e5072b06d104c50933019df8;
// music[6794] = 256'h4eff7bf594e864f418f979f4cdf65cef8debcbfcfe0154f5cdf6d102390d4c10;
// music[6795] = 256'h2a09eb070509bb064707c60317ff37faf1f503f31cee31f65dfb39f383f975f6;
// music[6796] = 256'h2fe726f269fd67fe430ab00ada0146058002f6fa6702ef080008190d170e6d05;
// music[6797] = 256'he703990cec12551328149419a11e0d1f981ed11b1f1a3f1daa1cd226823ff74a;
// music[6798] = 256'h4049ee45e142da44384ad34e31514653ad4f824a674afe489751a35907533953;
// music[6799] = 256'h13554e4efe3d5a31613cd9403f3d8541363557292031b138583a0b3bc2382233;
// music[6800] = 256'h24393944dc4394433645b24794497d442d454d48c942c237182fef339f398c3c;
// music[6801] = 256'hc8443b449742ff438e3fe04211497a491447f2407b3f4540333de0399d369637;
// music[6802] = 256'h224086495c492d3f5b311c2ad42c5b2e68343c3d563ccc3a2c36a6320741fe52;
// music[6803] = 256'h4752d641233c4a48265380548551724df147eb447c457a49184a08430947f149;
// music[6804] = 256'hcf469a48b13604295728c916501abd2bee2ba236c33e2434e229441b360fca18;
// music[6805] = 256'h6225ba234122e02478236d220c1e260c3e01d906e407f5064306220028fc2bfc;
// music[6806] = 256'hd9fe49f805efc7f2c3f419f0a4e973ecebf509f546fbc0ffccf41fefdae837ea;
// music[6807] = 256'hbaf60cf812f7c9f2ade7ebe335db06d24bd7fbda7ae067e4f6d95be0cbf31af6;
// music[6808] = 256'h98f1a6ef38eeb8e659e29be94ee806e410e1d0d770d5b8d9a6df9ee37fe4c9e5;
// music[6809] = 256'h7fd95bc572becdc013c357c4d9bf79b7bfb721bcedbbf6be43c417c2a3bf9ac3;
// music[6810] = 256'h55bcdbb8b8c7fac23ababbbc5bb373b847c1c1bef4c4a5bea3b763bc53bba3bc;
// music[6811] = 256'ha1b993b88cc281c49ac325c200baf0b5efb9c6bef4bf5cbdc6ba4ebf23c3c5bb;
// music[6812] = 256'h56b54bba85c651d044d4ecd45cd353d3a6d0a2c741c508d174e001eb8def3aee;
// music[6813] = 256'h2eef39f23cf053eaf5e5abea4aeba8e940f3ecef9be97ff02cefe1ed05e8d1d8;
// music[6814] = 256'h01d8ddd79ad32fdd1ee4cfe585e92fe1d3dcd6e293dfd4df19e32ee4f6e640e5;
// music[6815] = 256'h67e9f9e412da81e339e6ffe5a6f1eff037ec55ebe8e983e930e349e28aea4eed;
// music[6816] = 256'h8ef0d2f4e8ece3e618ec38ef60ede8e474dd31e01de545ec05f1acee52edfaee;
// music[6817] = 256'habf149f015ee66e686d853e161ef82edf7fd370fe00334fead08700b4409200c;
// music[6818] = 256'hae05fcfbc1018403ee00e507150e8d12f80842feca07a2ffb6edc0ef1fec4fe5;
// music[6819] = 256'h97e4c7e497edaef3d3ef88e845e344e92eeeb4e821eb8df209efd8eb0eef27f1;
// music[6820] = 256'h23f5ddf4c6ed97ed9def4aecf5ecc8f532fb6ef4c2f010f354f15af539f8d9f3;
// music[6821] = 256'hc6ef70ec47f16feecde519f12cf713f344f288ea51ee0bffc104390249032e06;
// music[6822] = 256'h56032906190fee120620bc2da1253a18361683199e1acc199921372d43288c1d;
// music[6823] = 256'h541d32212029cb29b321d820b116ec031b00dc023301adfc4b02b7101e0fb908;
// music[6824] = 256'hce085803c9005bfd98f81f00e704c7031c0ac60f440a0801d60020031c031107;
// music[6825] = 256'hb00431fc51ff6a0b1211530bb502a703240bd10be40796055001a7009b055605;
// music[6826] = 256'hb103a4051d01e9f77ef798fc31f4cfe970f544fddff5a6f78700a909e8074d05;
// music[6827] = 256'h2618281f66171c1d4221c61f0e1dc41c3b25fb226f1694153c17cd136f13080f;
// music[6828] = 256'h7011811544fcfbe5ddebeaf44cf767f160f48eff5ffefef9a6f357eca9f27600;
// music[6829] = 256'h3308000a4a0c870ec70b350089fc4a090411e30f251329194e176b16e31b9718;
// music[6830] = 256'h0d19241c371d0024601d8e185f21b32232215d200d249d2819282c27a1250122;
// music[6831] = 256'hde1baf1f1d23531fe0251b28382af82c6629e23217381434fa37c042304d2e4f;
// music[6832] = 256'h1650db496d41873f4638643a8f3e603be73e43432c40452c4a1b651e2f1f4421;
// music[6833] = 256'he1277a2d013093224f17a01c6d1e7e1db920d320d121de240324aa2888320d2d;
// music[6834] = 256'hce1d1f1b771d6722fd29e623ec19cf12f311461d461c2c16701a1320b624e51c;
// music[6835] = 256'h7516bf1a83179e16fa16f710de0eb01214155e0ce0038f0a4112750cf103090d;
// music[6836] = 256'h69199714ca17f626c6262f267b280920192028235b220725bb2026236524b017;
// music[6837] = 256'hd5192f2238243527f318bb03bd0143034ffec60330072efd01ffbd05bafd3df4;
// music[6838] = 256'hcdf0bffb1c0f930f810549006cfc74fd9dfcd4f352f16ffe460740fe0bfbdc00;
// music[6839] = 256'hfbfdcff81bf8b5f63af425fb8dfd1df675f840f1c0ea81f39ded70eedbf390e9;
// music[6840] = 256'hf9e60be381dce6dd45dda9dae6d9cdd648c92cceeee634e6bde01ee352d9b3d8;
// music[6841] = 256'hc8dd58d9e1da98dc6cd7abda7fe055dee2dd83dfb2e1bbde46cb73b6d2afe8af;
// music[6842] = 256'hb0b496bb80bdd2bfc9c26bc2ddbdacb4a1b6e9bb3cbac9bff9be4fbfbdcac8c6;
// music[6843] = 256'h11c023c036c04cc794ccc7cf8ad955e1f0e015e258e3a5dcbadabcdca5e253eb;
// music[6844] = 256'h4ae85be781e5c4dcbae2b4e861e4ade2dde4ceeb0ced64ea19eee9e962e670e7;
// music[6845] = 256'h3ee36cf7700f0f0b740ac70276f9e4004df90ffcde092603bd0583072cfb3cfe;
// music[6846] = 256'hdb09c20701fc03f4a6ecb7ebd7f31ff344f289f3bfeb96e922ef98f562fdf0fd;
// music[6847] = 256'h92f443e8dde292eb51f4f0f182f130f5a8f4bff11ff13af96f033503d2fc96fa;
// music[6848] = 256'h07fe8dff03024d06f5fea9f79cfef405f402eef947fb760001f319ea3bf0d9e8;
// music[6849] = 256'hf2e1f9e8c7e72ee5ceea88ed6af4c903670e100fc20c210b7f054b03d006d602;
// music[6850] = 256'hc1024a0bf50b820650fe93faecffc701c3ff66fa6bf3f0f30af383e961e333e8;
// music[6851] = 256'h2feecdee1ded03ed94ef96ec3feb23ef21e85de314e7b2e7e5e8eee62ee5fee7;
// music[6852] = 256'h8de86de926ea74e9e9ea5ff218f653ef03ee58efb3ed9bee13ed3be9ffe05ae3;
// music[6853] = 256'h77f2f4ec6ae3cfec31f4cdf19dea17e844efc5f4b2f09cedc1f91309250c1e05;
// music[6854] = 256'h2e019b07130e70108f0891fc11fc72f863fba809d7059c007705a0fa61e7a3e3;
// music[6855] = 256'hdeebbff27bf577f121ed0ded10ea97e987e9ece54ae9d6f16af235ea06e4cee0;
// music[6856] = 256'hdee216e8a6e845f01bf16de8adeae6e8dbedaefa99f319e9e6e48ae9eaf060ec;
// music[6857] = 256'h75ef94f136eafef318fb10eb72e140e428e67aed65ef0ded86f316f2f1f453f8;
// music[6858] = 256'he6edc8fc0d13320e900363fd9b015703ecfea2039f01fdf9f2f8eaf746f87dfe;
// music[6859] = 256'h4708d10a85fff2ec97e8c5edcbe6a5e994f496f516fef4069909050d680fad0f;
// music[6860] = 256'h99082905b004b5fe9efce1fb0efe3eff52f7dff3cff384f2c3f673fb43f8caf6;
// music[6861] = 256'h580145057efd8efc3bfc3afff80af10a3309b4105710fa100a12320bdc0f891d;
// music[6862] = 256'h0d202519b61b79241a1e121d9231694181401f3fa644c2442e42423e063a2f44;
// music[6863] = 256'h4f44613a9c4371484c44e548c441512f382d8f2ca723782db33567302d30db2b;
// music[6864] = 256'h15310f3a223477319f2e522b342a4028eb2ab5294f2e1c32e329272b8a2c7e2e;
// music[6865] = 256'hbd3c253e673c85475745673c7b411441433b4941194a05525658934fca3fd740;
// music[6866] = 256'h73486a41ec3a723c5d409d473a47d9427b41893c5f435c58c95efb564f56b158;
// music[6867] = 256'h4b57b253074e3b4c485187553d4c4c449c4d304e954f53555d3a21273430e729;
// music[6868] = 256'h9929c73635332c291e260d2e7f3035241427bc2e012a602b9727551c391b1c1b;
// music[6869] = 256'hc619651c501b1717cf15fa120c11731a34256a21331824180d1963143b16901c;
// music[6870] = 256'h681bda1589158016f1155719b912c3070409630672042301cff210f0a7f7ad06;
// music[6871] = 256'h7518e919b215360e310ce814780e110c9a16df174f1ccc1b4914eb107f04da01;
// music[6872] = 256'hc4ff0aecb9ec58f0f0e2d8e152e4e0e368e4c1dec7d829d6cdd51dd435d0c0cd;
// music[6873] = 256'h62cf56d189cdf5ce81d491ce8ac155bf03c8d8c361bbb4c08abfa2bb4cc3a5c5;
// music[6874] = 256'hb6c19fc62eca1ac61cc326be15bc6cbb55b8e1bd46bebfbb6ac15fc1f3bd89b7;
// music[6875] = 256'h1cb1b8b281b37eb80fc700d563d8c8d736d855d3cdd448dc2cdd34d952d2dad2;
// music[6876] = 256'hfed4ecd4d4de01e1b3d543c9a8bf07c2cbc262bff8c43ac466c0fcc357c503c5;
// music[6877] = 256'hf0c5bacaecc7b9bed4c8eed110c984c83ecdefc678c1fac91acf0ec8c8c773cc;
// music[6878] = 256'hcdce54d1aacfadd1add62dd03dccf2d3f9d399d5cbda92d390d30edb42ddfbde;
// music[6879] = 256'hf9d9f8d6d8db00dfc7d9e8d66ee3d0e414df88eddefd0a0228fd71fb6aff6102;
// music[6880] = 256'hc20634059605be02b6f5d7f486f88df852fb5afab4ecd0d79ed760e03ae253e5;
// music[6881] = 256'h51e0e8dfd5e4efe3f1e6f8e44be37de577e4f1eaf5f07de983de4fdf67e58ae7;
// music[6882] = 256'h5debf1e8b2e7ddec9be632e1aee5d9e68de237e5d8f214f30bebb9eefbf020f7;
// music[6883] = 256'ha4fa51ed35eb1ef2d6ef9ff059f353f22bee44eb01ef1df020eeccf001fe1c11;
// music[6884] = 256'hfc12de09c7099e0a1c0808082209a80555033a071708a008c107e3057509a4fc;
// music[6885] = 256'hbee8e9eb40f071ec8aef96f244f21cf0b0eef2f313f430ee02f13af14aeb6aec;
// music[6886] = 256'he1ea99e708eb29ecf9ed95eeafec04f10bebd2e4b0fa860e580ef30cf005f200;
// music[6887] = 256'ha508d30af30827096c02f9019d088e04e103cf0b000885fd3bfc8302ec06c707;
// music[6888] = 256'hae086204a3030d155423212268246426a0228725c025111f181f381f0718f416;
// music[6889] = 256'h3e22e927f021f9198607effa5f02ea007c02990d2a088a09b90c31fc53fa9502;
// music[6890] = 256'h6400ee03d507f408390cc308cb059e06a20350ff93fb4afa4efb7ffd54ffbafd;
// music[6891] = 256'h84fa76f531f401f9d8fcb0004203120723072dfc47f92f03920ab301dff65006;
// music[6892] = 256'hc10fa30140feed033a0a350c8a03b807331c91245720ec20f51ffa16e1112313;
// music[6893] = 256'h5d0e0f044607800ce906a50b8e11c60daf0ad6fb7cee26f6fdf8f8f35cfac800;
// music[6894] = 256'hf1040307e9fff1ffb4023b020f0be10d900a160b860d2e16d719db18f01c291d;
// music[6895] = 256'hc61c3b1f5919ce12ca19491fc01fce289230dd2fb52abe27312c8c30fa2eb72c;
// music[6896] = 256'he0305330232c2730862f9a30ab32922fe5327c2f352e533263325e45d850af47;
// music[6897] = 256'h6149fb48f8411544fc49984a8a4783445f3ef43df63eff3a6941de40f72d5323;
// music[6898] = 256'h7420db1b4d1c431f1d1e081cf91f0824f422a22391200d1b11206124c1223722;
// music[6899] = 256'h461a7113cb18c819d7153e18bb1725162e1bc2197915cb1c5c23821e7f16d513;
// music[6900] = 256'h44144e120e16d91c0e183b17111fbe190b12b811270f151195138711c9125e14;
// music[6901] = 256'hbf14b61a83265d2c532e9d315e2ad626b02d862cf8261024d526d824691fa725;
// music[6902] = 256'hd428172e502c6811c506fa08c6ffeefec2030a05a403cbfe9cfc2fffa9017707;
// music[6903] = 256'h1211810a09029e0417fba2f1bbf141f227f3d5efcff01df410f617f779f348f6;
// music[6904] = 256'h18fa2bfe800468ff25f8f7f097eb2df01bf008ec22eda0eee8edbaebd0e822e5;
// music[6905] = 256'h0fe198dbffd34ed344d9b5d6ebdc97f2a2f0b0e9a5f1e4e8e3e1c8e8f3e6bee2;
// music[6906] = 256'hf7e100e134de4fdeaddfdbdb69d9a9d49cc825bf4fbfe4c011bb2dbcbbc1a3bc;
// music[6907] = 256'h00b9ecbc05bfabbce1b7abb5d5b988bdc6bbeebdd5c5abcbafc640bb42be16c8;
// music[6908] = 256'h44c43dc053c23ebfa0c71dde37e39adea3e0c1e18fe343e022db65da3adbe3e3;
// music[6909] = 256'h60e7a6e026dc37dd53e2cae0a1e1aae8e9e802e77fe4a1efcc04f904b8ff9903;
// music[6910] = 256'h5106cd0a7b0bc102befaa5f92cfdc0037505c3fecf00410728fe21ef84e7aae6;
// music[6911] = 256'h85eabdecf8eae3ed26f1a4ea85ead3f144ec39e889f12ef400efd4f009f589f6;
// music[6912] = 256'h60f823f6f4f2c2f1b8efe9f2b2f6a9f9f9fc48f740f443f900f87ef4b9f6c1f7;
// music[6913] = 256'h3ff555f916fc0cfa2bff02fdd0f8c6011a03ef00a3035ff73fe600e5a1e5bfe7;
// music[6914] = 256'h7ef82b033606290dbf0adc07f60857073b096805c9fdfefdd80166057805de02;
// music[6915] = 256'h820021f7e0e734e4c0ec65f35cf2c2e84de54beac5e867e5d2e598e62fe6a9e9;
// music[6916] = 256'hf8ecb9e4cae196e525e5d2e829e82fe203e1a3e2f0e726eb09eb53eec3efdde8;
// music[6917] = 256'h7ae437eadaf0f4f1b2ef92ef58ee22ed56f133f29ff43df4fef0a8f84bf568eb;
// music[6918] = 256'h20ebebec40f4daf0f7efb4024108e4046309950c410c250ba409c307dd084105;
// music[6919] = 256'h5dff59035804b2018304ee01adf1fee2fae4afeca7f026ee4ae56ae1a1e112e4;
// music[6920] = 256'ha6e8a1e801e684e323e156e4e0ec44ed9fe700e94ae6b3e0e5e1e1e287eac2f1;
// music[6921] = 256'h82eb86e9c1eb3ee888e810ecb1eb30e770e6bdebf9ea87ebabf0a2ec9deb53ef;
// music[6922] = 256'hd5ed88f053f019e9c6e64ae778e8fbead0eadcf01205a011b30e4e0e320bb505;
// music[6923] = 256'h8806800543019dfecc06070b50026d06ad062801e403c6eca4d6d7dc5be09be5;
// music[6924] = 256'h64ea65ea2ff005f389f064eac6ef3cfff1029b04c402b501950def0f020a3708;
// music[6925] = 256'hb40432053108b50407feacfac8fa21ffe9fe86f6dcf74efcf2fae6fd2dfee0fa;
// music[6926] = 256'h38faef005b08f0044608bf0bd4049808140dbe0ddf130c15381309102c14c827;
// music[6927] = 256'h07341436893915359a320b384d3574365e40b4404a3e063d08362934433f4141;
// music[6928] = 256'h70307f2c642faa28bf2e0030d529df330b33972610250b27622a572f9b324634;
// music[6929] = 256'h74369a379f34dd327f3329344b31b32d6b2f2c305430c5329933be312e345441;
// music[6930] = 256'h8447e0473d4eae4e68500d539b518452ea4a77463149c345034600483248a444;
// music[6931] = 256'h27410e478f46d54a9f5bee5a5454bc570459765816562a54e5538750174f594e;
// music[6932] = 256'hfc4c764c6a4db755ce4f1238c6313b31532a302d9e30c42dbe268126472d362b;
// music[6933] = 256'hd82a2d29c025f728f0248327602c25235c22be259f248b22961de91d031dfa1b;
// music[6934] = 256'h892281246b21652250276328ac237a219621f01fc41f4522931f6819961efe25;
// music[6935] = 256'h3a1d1e14b31647186915730b7a008f06df161d220a22101c0115830ca9101714;
// music[6936] = 256'h500aab095e0c500eda11fb10e3134b14bd11490a7ff7dcf078f3f9ef0aed35ea;
// music[6937] = 256'h81e81ee557df36e024e10cdec2da2bd4ebd184d65ed30acf67d246d1d7cb10c9;
// music[6938] = 256'h3bc56cc42bca71ca23c62ac71acaa9cb64c4eabfb4c632c32bc1f7c463c33ec5;
// music[6939] = 256'h2cbc9ab99fc5c2be28befdc574bc3cba92ba9ab26ab81dbdfab8b0c7fdd572d0;
// music[6940] = 256'h76d0dad123cf4ad2f0d34fd570d337cc03ccd0d05ed38cd266d5c9d91dcd27ba;
// music[6941] = 256'h3cb957bfd7c05bc295c26ec3f0c2fdbcd4bba6c1e3c48ec011bea3c2afc5b9c9;
// music[6942] = 256'h11c8dfbf87c448ca54cafdcc6ccc58cf77d05bcbb7cfd4d081cd16d545d580ce;
// music[6943] = 256'h12d078d211d984df87deebdc27d7b5d31dd6f4d83cddf8d74ed2f4d851dec7dd;
// music[6944] = 256'h27d862d788e69ff408f506f4bef51cf407f6e3f8e8f74bfac3fac3fadaf94ff5;
// music[6945] = 256'h09f6b6f514f591f16ee3dcdd5ee251e50de5a1e31be4f1e0f1e0c7e5ede4b3e1;
// music[6946] = 256'hd9de81e29be6a5e11ce08fe4c8e74ee5a7e267e5a4e2f4e37fedf5ec2ceb44ed;
// music[6947] = 256'h77e95fead7f270f659f652f451f0b3f1def0d2eeb9f70efa4af570f869f920f9;
// music[6948] = 256'h09f47de971edadf40cf491f226f24dfff50e6a0d0507a406ee0833079803a802;
// music[6949] = 256'h4b0471086408470bc40c09031e050f060bf5d3ed81ef08ec49e795e7f1eb29ec;
// music[6950] = 256'h7feb46ec75f071f1e8ea31ed1ef0aced25ef3cecf4ea6bed03ed81edb1ee58f1;
// music[6951] = 256'h8af393f5e2f298eb9ef2fdf83ff14bf12bf42ff6f6046d10830f3e103d121f11;
// music[6952] = 256'hc20f28113b133010f10d030f870cb9084e09ae09c302c808fe1ec3245c23ba25;
// music[6953] = 256'haa2114244422f6193c207c223f1b241fe8259c257c26032b46251e0ffd01d006;
// music[6954] = 256'hbb04d40039078f073a0120ffd20067017ffe8800f1040efdaef405fb4dff5bfd;
// music[6955] = 256'hfefd05fcf3001209ed03e0ff0b0138017502b8fe0efcd3048809deff67fc9c02;
// music[6956] = 256'h8402adfe80f95ff938fbe8f92c025e03edfc6505ae0e020c68fd52fcad0e110c;
// music[6957] = 256'h7906b414e71fe523fb2020200021791931178518b9171a137d0c94110b11350a;
// music[6958] = 256'h5011970d93fd7df927f7b8f55dfa33f9d7f7d7fbb6fa6bf7c7f9b600a7047c02;
// music[6959] = 256'h640190ffcdfefe01a403720a7d10b413661abc163b113c140617eb1b5b1f0322;
// music[6960] = 256'h22240c235b25d827c029602e6e2f2f2d212ff82efe26dc272e2e6a2bcf296631;
// music[6961] = 256'hae34242bf42d96341f2c4938c8485846f647e7456545f54670429f44c044b343;
// music[6962] = 256'h0f43f63d0041fb448446434aed3e5425e31dfa26e023271e6b2072205d20381f;
// music[6963] = 256'h941f2728222c59224a1cb01fe720eb20041f6a1ca61cd11d10238e232f200e20;
// music[6964] = 256'h481f7821d620721f6b21921c2f1da722c11e4a1a6b1bbe217225991e251ab31f;
// music[6965] = 256'hfe221c1c5d163b1afb1b1519ba19ec1865155a125d19062a6829cf252530be2c;
// music[6966] = 256'h6027282a1125b7210c211b22ff28072b31247a219424c018cf0805097c0d6710;
// music[6967] = 256'h520cda06f9072c0434006000920223041fffd1feab0048fe50fd66fc7203ad0a;
// music[6968] = 256'ha30296fcd2fe47fbe1f553f7d7f65bf185f591fff2fd24fbaafd76fc6901af02;
// music[6969] = 256'h29fa3ffe4aff2ffb82fd69f45ef2b8f7fff18bf20af133ec37eb09e04dddeaef;
// music[6970] = 256'h60fe9df845f0faf022ef76ea33e6bfe70aed2ce9d1e44ae58feab3eb8be3e2e3;
// music[6971] = 256'h02dec1cb37c298c08fc43ec2a3bc60c09bc0a9bde6bd97bfeebc88bb38c0b3bd;
// music[6972] = 256'hb4bea6c02db9b7b86db81dbb62c0c3bd0ebe59bc4abd6dc333c2e2c24fc704cc;
// music[6973] = 256'ha9cd0dcef4cf45d103dc34e127da3dde2ee537e323defbdb35de79e224e68ae3;
// music[6974] = 256'hffe182e0c3db62df7aeaddf9b0fdd2f6bbfe2c0153f889f9a8fcbefdfefa55fb;
// music[6975] = 256'h3206d6047cfd830481047cf35ee7b5e60ae732e88bec1deb4ae8ddeb78e986e5;
// music[6976] = 256'hcfe90fe9a4e559e774e761e7c5e988ea5aea65ef6ef432f1f0effaf191f294f7;
// music[6977] = 256'h01f8cbf47cf8d1f626f629fcb4f82ef654f875f9c1fe74fdb9fcc9fe70f7a9f3;
// music[6978] = 256'h78f35df7bffcd2f777f971fd67fb29fae4fa4b0c3115ba03e6fcc401c3019eff;
// music[6979] = 256'h8401c905b70091fede0575089a056f0387064502d0f02fea07ec82e720e910ee;
// music[6980] = 256'h54e93fe32be164e486e775e5f7e7ffe78fe3bbe596e645e7d7e8b4e765e56be1;
// music[6981] = 256'hb3e4ebe9d5ebd4ee63e9cce30ce9bdee08eed0f0f4f456eccbea30f3f7f442f7;
// music[6982] = 256'hbbf483f214f30ff06cf43ef50ef290f260f25af2e0ee0bedafe9d7ed7eff7d00;
// music[6983] = 256'h7a00c706d400f3007c0190fe8c029a0017fdce00000486002100b304fafcd7ec;
// music[6984] = 256'hdce3cae6d6eda1ec3dea11ebfee8abe648e59ae3e3e29de415e921ebfee78ce5;
// music[6985] = 256'h00e6e5e505e2b3df26e60ae800e452e7fae7b1e82cef49ee73ed61f32ff47bf0;
// music[6986] = 256'h72f2e6f2c9eaf9e900f2f9f5cef5b3f5a9f30ceff0ef6bf079ef95f31def86ee;
// music[6987] = 256'hecf38eefcbf43ffc21fa35faf6fa4003680a8a09150ded109111170cdb066d09;
// music[6988] = 256'h8f083103210060ff78f5e0e9b0ed1ee9dddd36e243e867e795e2dfe018e2bce3;
// music[6989] = 256'h65ed2bf49df315ece9e671f56bfa39f4c7fe9107f4094e0c63090c055e014a03;
// music[6990] = 256'h2f03e100e504450102fd3e007efea9ff9a019cfc3efb52fd2b00af0092fd7502;
// music[6991] = 256'h080535fe6b011d0563028506e6051b0bc3204727d12248276e2aa82ac52c7c30;
// music[6992] = 256'h2931712fc631b0333d36be37933619396031ce225922dc273628672485241628;
// music[6993] = 256'h49254425fe2bde2d7d29f227e32c5233c636d2361d390038d531dd333233d033;
// music[6994] = 256'h133ad434743482385b38813bb73566339135b5328c3833393e341339e043b14e;
// music[6995] = 256'hf94ccd458a4401443346a747d746ad45ac42cf458846213da64375545353204f;
// music[6996] = 256'hc950a54f0252bc5783588554d2551254f94dd852d452a550b4521444fa345f2f;
// music[6997] = 256'hdd2dd6315f30bb2f6b31862fac2e382ac328ab2b062afe272025ed217e24d629;
// music[6998] = 256'h282de52a192688236e20c8216829802c3429b1238e246425811c831b61232427;
// music[6999] = 256'h2c267f259d28fa21661d51249d25b525e2233124c7239b19b619411a07194b1b;
// music[7000] = 256'hee15a41fce2aea279e284a22051d691c0a15d410950efc0d190e9f0c270c2007;
// music[7001] = 256'h4c04800505fd79f559f7fff3b1f1e9f5d2f11bf04ff6f8f504f130ee4fee43ec;
// music[7002] = 256'hffe7b3e659e52be48be16ce0d7e1e2d987d22cd60fd471cdb3ce9acb9dc484cc;
// music[7003] = 256'h2bd47dcefcccedca19c56ec93dc98fc326c8b9c828c6b6c6d3bf94bdd8c018c0;
// music[7004] = 256'h1bc24ec21ebf0ebed2bad8bc4dcd2cd9f6d7fcd801d403ceffd243d226d28ed5;
// music[7005] = 256'hf5d1b5d0ddd452d9a0d52dd5c3d8c3cae0bdd2b8beb895c0b8bb5ebc2bc2f9b6;
// music[7006] = 256'h35b802c282c015bd86bc69c04cbfc1bdb8c449c567c0bcc148c61dc5abc059c0;
// music[7007] = 256'ha0c1e8c35cc781c9dec7c7c6ccce64d4ced247d5abd64ad3ecce0ece27d527db;
// music[7008] = 256'h7cd903d714d588d46ed8d1d6b8d36cda7dd9f8d50ee0bbe967ed58ebc2ec31f4;
// music[7009] = 256'h08f166f11af7f3f1aced21f072f579f655f2f3f20cf955f8b7e634ddc9e0d9da;
// music[7010] = 256'h7ddbe8df60e1bfe619e1c4dc39dff4dcf9dd5fe2cce768e546e2c3e71de77ae8;
// music[7011] = 256'h2ceea4edc3ebaee87de7bde8f0ead1ea84e72feccdf246f230f060f13df0d6e9;
// music[7012] = 256'h5eebcaf033f247f308f194f215f658f607f4a6f0a5f426f2ddeaf6ed82edd0f3;
// music[7013] = 256'hd706590ec1078603c706a606a4063d09f804650317069b06df063605d402c402;
// music[7014] = 256'haffe04efd8e708ed44e621e603f1c9ed55e990e9b8e92ced29ebc5e7dfede5f2;
// music[7015] = 256'h51f0a9ef43f236f5c3f5bfefd1ee20f41cf318f1fef0f0ed18efcbf6c3f94bf6;
// music[7016] = 256'h41f57cf707f9a1f661f484f94afe55f9cffa5408820aed06c40b980de60cf20a;
// music[7017] = 256'hc409990a2f071e069c0fe821fc26b11d951e921e8e1b231ce11c611da417fe1a;
// music[7018] = 256'h5a1f4e1beb1e911a2219a618d90270fa5a01c1001000a6ff33ff4c02c9044901;
// music[7019] = 256'hb4010106da0212029c00d6fc9601c802b0ff1201c5fc4afaddfec2f975f91f06;
// music[7020] = 256'hbd063e041c0c9a0fa408f402120371021a016ffe8b0193079c04a505a702b4fc;
// music[7021] = 256'h15fc51f503f763f945f610fa06fb0c00d8061914951d1317fe1f1a25e623052c;
// music[7022] = 256'hb4231d220724be1dd81ffc194e18a21ae913da145a0ff6fd64f4eef18aeeb4f0;
// music[7023] = 256'h76f610f2e2ee8df0bbf2bdfbd8fc18f78bf941fd82ffa600ff03960974071107;
// music[7024] = 256'hd70a9309d10c450e0c0b880de410ee19771ebf18541c951ebf1d4f21d6227b26;
// music[7025] = 256'h1e262225022a842b922be52a8f2c412c64267329b62d332b422b522cbe35c945;
// music[7026] = 256'h0a492b474049e3451543ce43ca42e24096411d46a144ff425c46ad4363430a3b;
// music[7027] = 256'hc426c32147257c25f8266e28bc27e42403276d277a241427cb254b2254238f22;
// music[7028] = 256'h96227326b3267121f22078223b1f4b1f852154210a20871f1222b621311f6d1e;
// music[7029] = 256'h471c5d1d1221eb22b7226e1e261d4f1fa71d921d7d216122901cf919cf1c8c1a;
// music[7030] = 256'hdd19dc171718ee29c534823363337b2dd62ddd2c5b23ee235f27be28d626c723;
// music[7031] = 256'hc1277e24b221e123f715c1070e057502d6026a0686081b07b106d1092809ee07;
// music[7032] = 256'h9407070656077105e700cc00510310060a06ee04a00002fa8dfe11075a070606;
// music[7033] = 256'hd804bc02ae014cffb9fb79fb29fcedf9a4f832fb95fda8fa29fbb701b2fe82fb;
// music[7034] = 256'h7cfe34f941f6daf72af5def459f17ef2780245081c013a0045009dfbc2f591f1;
// music[7035] = 256'haceff0ed15eedfeb04e88ce9d6e757e586e4d6d5f1c7e3c962c7b4c2bfc748c8;
// music[7036] = 256'hefc3abc2d1c1dfc352c50ac4c6c2e6bf03bf43bfe0bfe8c27fc2a1bf76bf01c1;
// music[7037] = 256'h5fbe0db947b85fb8aeb88bbd48c35ac3b8c07bc4b6c615c4e0c4c9c603c837c6;
// music[7038] = 256'hc3c5ecc75bc628d0aae0ade03edb6add1ee0a4de67dc81dc17e36ef0aef75df8;
// music[7039] = 256'hecf946f9cafa02fd5bfa5df80df777f961fd0afa2ff849f893f94dfb1aec68de;
// music[7040] = 256'he2e2a3e4c5e587e85be9b6ece4ebe8e97ee9daea8fed6be997e821ec76ea6ceb;
// music[7041] = 256'h38eff0ed58ea69ebd2ec7aecf1ee57eec2ed7df0a0f334f64cf544f862f986f4;
// music[7042] = 256'h63f579f684f77bf6ebf3c3f785f639f710fccffb87fe86fbeef559f85efbaafb;
// music[7043] = 256'h16f8d600721174139911b2122f14a914611355114c04faf8c0f91efa11fd7bfd;
// music[7044] = 256'hbff9bffe22fb69e7c4ded6e120e4d2e849e8e1e698ebfbea7aea46ec50ed48ef;
// music[7045] = 256'ha6ecc7ecd6eddaea16eccdebafe97be976ebb6ee21eb18e847ea50e932e864e9;
// music[7046] = 256'hfaecbaf079ef0eee59ef1beedcec1eedc4ee42f217f040ef09f280edd2ee77f1;
// music[7047] = 256'h67ecb4edd0ed0af00ff593ee61f54d080b09d204000831084d04bc038b077706;
// music[7048] = 256'h8b0243016afe22013a044cff08024ffe60eb87e511e66fe4c4ea49edcfe9c0e7;
// music[7049] = 256'hc7e6ace8b8e848e51ce79eead4e825e9dbe9f9e83eece8ea76e740ea47ea81e7;
// music[7050] = 256'hc4e6b1e7e4e770e600ebbef05feeaeed50efbcec8eecc4ee74ef6deff7ef63f2;
// music[7051] = 256'ha4f0d9ed2ced78ec58f228f30fedb8eeffefb8ee08efb6f9c90a360b3a07e109;
// music[7052] = 256'h3f080101fffad801e90475000507d00b330a8d069c03cd06b4ffa2ee22e878e9;
// music[7053] = 256'hf9e5a7e86ff23cee57ea15ec57e447e025df62de52e19ce0d8e346e787e996f3;
// music[7054] = 256'hf7f816f3bdead9eac5f199f5ccfcbf033305e10b880f570ab509210bb7078703;
// music[7055] = 256'hdcffa3fd79fc4cf92bf813fa22f9c3f9a1fc54fa23fb99fe4afdac012f041901;
// music[7056] = 256'hc70d101e29202c225026c72558265e29c72ad72b172f3431772e7f2b012c0f30;
// music[7057] = 256'h3134392af21a7d1a6e1e0722cd25fa2507295f27dd23b4262629172daa2b7a29;
// music[7058] = 256'ha12d2f2bb12af62c2e2d9e31bc3038308c314a2d5b2d772fae300f30fb2e8a35;
// music[7059] = 256'h6c36da3107355236b633fa32c1313e33e936f33440336734e0304834ff3e0a44;
// music[7060] = 256'h0849fb491546f5439a421c4e725a6b561a57a75ad5568e57f756f5523954c657;
// music[7061] = 256'h4e5814540651564fd84e714f96434237f937b3371738613bb93bd5379a33ba35;
// music[7062] = 256'h7b34e13038334732b030193382335e300730aa2f7f2ba22da52c3626d3273c28;
// music[7063] = 256'ha329bf297b23ce25062bda2ac428b1279f267121ed223b265c22a620da1e091e;
// music[7064] = 256'h4e1fb41d891d86200726cd27da230f21901e4023ac313039b736ff33bd316e2e;
// music[7065] = 256'hdc2ce32d152d302cb52ca824321b5c18ab0f4e0c130f6bffc6ef42f06bf0daf3;
// music[7066] = 256'h6bf919f701f6daf605f5fef36df1f8efc3f14df1bcf1bdf17eec9fe9cfe949e6;
// music[7067] = 256'h55e3eee347e0d1dad0dcd2de56db8fd8add54ed50ed9b9d68cd39bd50bd31dd1;
// music[7068] = 256'h62d185cccccad6cbe8cae6c800c57dc43ac608c7b3c4bec2e6c5e8c09dc029d1;
// music[7069] = 256'h11d94cd9c8d70cd42cd61cd4bed292d5e8d4b3d6bed35ad199d425d17dd187d0;
// music[7070] = 256'h20c3ebb80cb7debafabde1bb85bc80bc36ba90bc8fbdcfbb03be91bef7bc70be;
// music[7071] = 256'h40bd30bc3fbf10bfafbc80bb77bc67bf60bf4ebeedbfa3c2adc4a8c4fac53bcb;
// music[7072] = 256'h4acdeac944c931cd46d0ebceedcb89cb44cc3ad08dd4abd344d3e2d417d838d8;
// music[7073] = 256'h8cd411d875d970dde8ee41f4ecee8bee84eeb1f292f280f056f72af770f22ff3;
// music[7074] = 256'he6f418f83ef736f658f354e4a1ddd0e1e2e034e25ae1addfa1e4bee262dfcbe0;
// music[7075] = 256'h7fdfdae167e339df9de0abe420e429e444e649e7e8e7cce621e4e7e5ade8e0e7;
// music[7076] = 256'h7ee721e61ee5bee839ed9aeec5ec1aec1eed4feb33e909ecc4efb7ecb2eb5aef;
// music[7077] = 256'hdeec67ec3cedf6ec30f15defeaed81ef86f40e06ff094e053b0b740ab9085108;
// music[7078] = 256'hd1050908d006970526060a05410626099c0835fc7bee6feb80ebf8eb11edf4ed;
// music[7079] = 256'h26eff3f0e1f0daef5bf1aaeeb1edeef15bf260f2f2ef2bed21f0c6ef13edf0ed;
// music[7080] = 256'hc9ee86ee78f2dff468f1b3f137f16eee65f028f14ef187f1c7f23ff7edf5d5f1;
// music[7081] = 256'h8ef371f4fef26ef2fcf320fa81faaff74c02480b170ab7052d049713d1213b22;
// music[7082] = 256'h8622001f5c1ec81ff11b9c1e0522ea1dcb19d51ac81e531e891c061dcf140806;
// music[7083] = 256'h1f03d406b806a0077206400462024a014e04e102eb00f8011b00f50041019dfe;
// music[7084] = 256'h830019042b00c3fa29febd0095019904bfffb0fad8fea2021d03c5083f0d9b0b;
// music[7085] = 256'h8a0d630d0e0bb00ce10ac307c002b6ffe904200abf099d03200161ffdef7fbf8;
// music[7086] = 256'hf7f9f6f8f00886179c151b18f01f73232227801e3d16802225252b25902ee827;
// music[7087] = 256'hff2086234223b218c804bcffdb023c0039ff8dfa77f784f69df2daf167f3b4f4;
// music[7088] = 256'h08f30df262f544f635f54cf5fbf700fbcefa0afa24fc170202058c036207860c;
// music[7089] = 256'hb20c010d700ee510b4157117bd17121a5d1a061eb42284203b1f2c20de24002a;
// music[7090] = 256'h54250b24fa25ba24f82aef295428483c1248e44301469c48b349f24902485447;
// music[7091] = 256'h0144b045d649604576454c49584c084f7d3ed32ab32ccc30ab2e9f2d072faa2e;
// music[7092] = 256'hf02a292de12c4629f12ba0282d25fa250a26152abe26e722fd2515234122ab23;
// music[7093] = 256'h0a24c926a02506241b241d232e22dd211622c01fc31f93246c25da20fb1dba1d;
// music[7094] = 256'h091d3c1d051c841ea4234820c91fef1f241c851faf1cf21ce82c83345332ad2f;
// music[7095] = 256'ha52c8c2cec2b7a2c562e492c5f2c102ecb29fd26d9270e2bd12af21a51105f13;
// music[7096] = 256'ha71130116f0f900d2c0fbf0a440b410ca808ed0bd70d9f0f0c11490cd60a000b;
// music[7097] = 256'h2b06f80388071407db053509ff07d605f4048e005ffef803be0c220a50026304;
// music[7098] = 256'h9a05f5fffefab0fab5fd93fc46f8eef8c1fc53feccfef0fe35fea9fd52fd40fb;
// music[7099] = 256'hb8fd370ba010ec08f4079507ee046104c300e2fd9bfaf7f9e4fa94f8d6f85ef4;
// music[7100] = 256'h16f2e7eea9dcc9d30cd328cebecf36cd9bc9d9cb6fc923c63bc544c41bc34dc2;
// music[7101] = 256'h4ec06dbdf4bf65bff2b82bbac3bc26bb0ebc81bb05bb32bfadbe78ba4dbd2bc0;
// music[7102] = 256'h01be6bbe4dbf12becfbe9dc2bbc530c4c8c3c6c5bdc58ac561c51ac837c8e9c3;
// music[7103] = 256'h18c743c6b3c6ead652dd28e18af10ef5e7f2a5f89af878f551f83efb9bf60bf5;
// music[7104] = 256'h7cfaf3f849f804fc71fb4afe22fbd6ed22e974e80fe614e786e725e6e3e407e5;
// music[7105] = 256'h35e50ee600e903e84ae669e7bae613e794e93eeb37ec43edf9eb3bea00ee89f0;
// music[7106] = 256'h18f084f0d5edafee55f219f2e6f171f08df0c2f23af4ecf793f678f349f7e2f9;
// music[7107] = 256'h2cf921f89ff740f94bfc74feacfc23fbdef9daf98506cd13bf14c71482156416;
// music[7108] = 256'hf71769146110c41022154016d81214186418e60b2307dcfeb0ef09ed51ecabe8;
// music[7109] = 256'h6de808e817e891e703e8e7e72ee65ae9e4e928e6d2e61fe727e5b0e4d9e5c9e6;
// music[7110] = 256'h3de862eb87ebc4eb24efb6efa6ef85efdbeeacf044ef1eeb40e9a2e871ea1fed;
// music[7111] = 256'h37ef4bf0d9ef4ff1c0f036ee58f15ff388effbed44ef7aee41ee09ee4aed29f6;
// music[7112] = 256'h5c021e05e703360174029707f105f00328042c03bf024002b905f6058903d608;
// music[7113] = 256'hd60240f2dfefcff0a3eaa5e81eea78eabfe846e7b9ea7eeda9ed01ed85ead2ec;
// music[7114] = 256'hbfec76e6b4e8bdedd4eb4eeafeec48ee00eae6e84fec77eb4fe942eb64ece1e8;
// music[7115] = 256'h6fe9f5ed6eec5fea0aeb8cea4feabfea7dec92ee7bef25f23bf3e1ee2eede8ed;
// music[7116] = 256'h21eee5f22cf056ec48fab105d705c305d905ea0705064c036104aa032c086c09;
// music[7117] = 256'h34ffa6fb08007d08390e23008bf29bf3e0f326f60ff4b7eed8ef61ebb8e7b9e7;
// music[7118] = 256'hd0e938ed00e684e40ee423dbf4dcfedc99dcdfe0cfdf92e4cce948eb7cf29ef8;
// music[7119] = 256'h97f019e6e6eff0f72bfb6c07d807ad09a910920a62073108d30749060803e103;
// music[7120] = 256'h13028dff4afec1fb9bfdfefce8f999f8c9fb8f0a5814c9137b15f9141118041f;
// music[7121] = 256'h621e661df01d892085263e28ba2a942ef6300d315723a4153d18261c9a1dc81f;
// music[7122] = 256'h2b1f3c20ee21961f781de320a9256123f21f7d233d27e528a92a8a29e329902c;
// music[7123] = 256'h532baa2b692e072dd72ca52e7c2f162f9a2b7f2cf62d6d29c42a2a2d472b3d2e;
// music[7124] = 256'h7831f73028312e311730f13386367f300330b5302630e2339a2e1d394f565b5d;
// music[7125] = 256'h585cae5fc95cc45aee594c5b575a9b58475bf1568755335b60588e58d959354a;
// music[7126] = 256'h2e3d5e3eb33cb33c0c3e8837ac3667397c37ae36b533fe3212342c2ffc2e8d32;
// music[7127] = 256'hfb30da30d030302df72ec632c12edd2da231892df329442a9928d72a562c5929;
// music[7128] = 256'h2d286f27ce2726298e284428a927e8254125de24c022322116217a2032207322;
// music[7129] = 256'h3924d51fd923d736b43ed03cf63bb237d1365433aa30e931bb2da82fa42f0230;
// music[7130] = 256'h82359f2f2f368e35c813e1041006cffd39fb07f8bff441f76bf76cf55df4a4f4;
// music[7131] = 256'ha0f4b5f320f36df309f53cf65ef7c3f63bf202ef3feedaebd9ea5eebf6e74ce4;
// music[7132] = 256'h7be610e7ace18de030e180debedd0cd860d343d557d2c7d0b0cf04ce25d3a6d3;
// music[7133] = 256'hb6d089cecaca1ac918c795c473c286ca84d902db3eda6cdaa6d472d48dd489d2;
// music[7134] = 256'h15d2b4cf95cf3ad2c0d714d9c5d369d61cd356c079b7fab9c6bcacbd27bab8b9;
// music[7135] = 256'h51b829b5ccb989ba16b6c7b4cfb5aeb986b878b681ba79bbaebb95bea5be08bc;
// music[7136] = 256'h62bceac0a0c2b2c1f1c1dbc082c094c3bdc531c886cb1aca00c91ac90bc780ca;
// music[7137] = 256'h48ce7ccdcdcd6bcfbfd369d531d1bcd07ad3cbd334d37fd4c0dd6aec2fef8eeb;
// music[7138] = 256'h5ceed5eee3ef62f0b6eaa1eb12ee66edd3f075f155ee60f194f6b4ec81dd8cdd;
// music[7139] = 256'hcadfbfde92df31dec2e095e15cdc6adeeadecfd8ced83ada6cdbcade0de092e2;
// music[7140] = 256'h10e315e252e306e339e588e784e719e6dfe16de3f2e5a3e319e337e316e44de7;
// music[7141] = 256'h79eaa5e80be7aee919e70fe756eb3fec60ef02f05bf088f276ee21ed20f198ef;
// music[7142] = 256'h54efe5feef0d300ac507700cfa0b180b0b0b1c085a0432076a0d6f0bd109f50a;
// music[7143] = 256'h45099e0888fef4f1bdf268f198eff1f1d7ed9fea4be90aeb9ced1ce908ecaeee;
// music[7144] = 256'h7be945ebbaeccdedf2f0faeed6ede3ecfcec55f0cff03aef47ed50ec7af08bf2;
// music[7145] = 256'hdced34ec82ed0deefeed3cea1bece3ef10eee8eecaed66edf0ee8aed94f1e2f4;
// music[7146] = 256'ha0f508f549f19ff2bff185f21100be113f1f4721551e331d961c34211d21981d;
// music[7147] = 256'ha71ffe1c261d0123531d0c1bc921e31599053b07f1071507980a35081d069e07;
// music[7148] = 256'h4405c902b303e40312031b04f204ca034502a703e40543031900f90092023c02;
// music[7149] = 256'hf9ff6a00d704b006f40301051409e7035ffc1ffe8303f10603071908180a3b08;
// music[7150] = 256'ha108b90afa0a540a4108940766031d03780b6b053e0102135d1a78137211ad11;
// music[7151] = 256'h1914c2164d18641c2921b1240325c01f9a17f219a2241223a11cec1a3814070e;
// music[7152] = 256'hea0b5f08b906a305affe66f9a7fbeaf762f19af2daf2eaf316f66ff4c1f30af3;
// music[7153] = 256'h71f54ff8caf7c4fa2afaa6f810ff2801a3fe3101eb05d207fb079709960c5f0f;
// music[7154] = 256'h431015103e122d150f14e3113d15561aa81bed1d36235f22f61f04255f241a2a;
// music[7155] = 256'h8c3e9641983e10456942c3419a47924a65499246cb4a1b4a40450748d046ce47;
// music[7156] = 256'h6d47a537c52d2830f82fa12e4d2d712b92298a2511250d28262741275828ce25;
// music[7157] = 256'h0f26632a912b522a122bc3281625d425d02427253b273525c725572727278426;
// music[7158] = 256'hbc2366223821e9207c22ae205120202360234222f91f421cc31e0e22371d921d;
// music[7159] = 256'h8921232011227e213a259e35c839e4334636c938fd358e326d35d63938351f30;
// music[7160] = 256'h272fdf2cd62b572cf32d022a991afa116414d013d3141a14f30da90cc30a0f08;
// music[7161] = 256'h8009a408bb08e009da07bf08800ddc0e830ab7091a0ee00e860c330af509fb09;
// music[7162] = 256'h3d08e50821084e055f04e9033304170234006e02ea05410af908060218feedfb;
// music[7163] = 256'h11f901f84cf94cf7c0f5f9f9a5fbe7fa0afc83030011d213d90f03123a136e10;
// music[7164] = 256'ha20dd90c290cf0098807f8031e016bfe96fcc5fce0f377e474deb4dcb3d7acd6;
// music[7165] = 256'hd3d6d0d1ffce64cf53cdbdcd1bd02bcc7bc83bc986c6e2c444c644c457c2ddc1;
// music[7166] = 256'h2dc2bcc16abf3ac077c082be08be4ebd1cbd2dbc1abb2dbc2dbc15bc50bc52bb;
// music[7167] = 256'h6dba69ba3aba65baf0bc1fbd93bbe2bd11bfe1beb8c0e1c3b0c576c58ecf20de;
// music[7168] = 256'h87dd18de32ecfef47cf4b5f40df756f8f8f6fef3f5f208f6bbf690f511f717ee;
// music[7169] = 256'h3fe03ae0cce106e021e16adf63dfc4e045df7de019e2dce385e53ce3c0e304e6;
// music[7170] = 256'hb4e41ee503e701e69de442e68be8a4e80ce97dea21eb5febb0eb36ecd2ed7def;
// music[7171] = 256'hb4efbcef3cefc7ee1cf089f0d7f08df1f7f1cbf446f5a2f3e7f5a9f9dafa16f9;
// music[7172] = 256'hd8faa7fcd6fc440a0217f61592166b186819ec199818761aea192d17c4149b12;
// music[7173] = 256'h9a15a2145e1384168b0be8fb61fbe8fdc8f550e96ee570e6c9e479e5e9e661e6;
// music[7174] = 256'ha5e72ee7e4e4bce5d2e69ae670e6c6e5c9e636e900ea54e93be8ece7c1e861e8;
// music[7175] = 256'h48e7bae81eeaf8e88ae99ceac2e82ce78ce6c3e68ee8c0e8a8e760e78be7fee8;
// music[7176] = 256'h1ae978e806ecf7ec23eabaebdeeb0eefedfe710969084609ca0a070b870a6409;
// music[7177] = 256'hac0bd00ce70a3c080706bb0754071c07a3067ff7cdeab5ebb8e937e968eb37ea;
// music[7178] = 256'h56e905e88be880e9f7e8c9e957e89ee73ee909e94bea98eb41e93be8ace997e9;
// music[7179] = 256'h4aea66ecd4ea39e86fe8f7e97bea1ae973e81be893e8f1e9fee8c2e962ea49e9;
// music[7180] = 256'hc7eac5e81be792e9e3e8ade808e9a6e959eba7eadeea8de9c3ef680094051406;
// music[7181] = 256'ha6089e056505d104eb04ff0624047c0550054b0176023d0271056004f8eed8de;
// music[7182] = 256'h96e3afe769e7f8eceeefcdedfdeef3f0e4f074f02bf0f7ee6bece1eab3ec93f2;
// music[7183] = 256'h71f200eb37e8b4e52ee27be16be07de253e646e885ea7dedd7f16df7daf691ec;
// music[7184] = 256'h4aeb6cf52efa59005f08260a130b9c0b350b6a0a580961065802b4013c02eaff;
// music[7185] = 256'h51fac0ffd7101715bb138e16d214d21346159c18011a6c189c1bac1ca41bbf1b;
// music[7186] = 256'hb71a891e591c3a0e46063f081e0a390b430f5311c00f3512af15ea1599178a18;
// music[7187] = 256'h8b18a11cae1e311e4d21ce2253238625ea240b26a129fe293e2a772bd72bff2c;
// music[7188] = 256'h112e702ed52faa3032306b30cf2f5a2f4330462f742f0f31ad2f602f8930292f;
// music[7189] = 256'h7e2e773071316c32e032f32dfe34124aa44d5a49c84bed4844509f5ea360be5e;
// music[7190] = 256'h4e5d2b5edf5ea55c655bf058025b6d58ec45863aaa3bd13a773a813b8c394938;
// music[7191] = 256'h0139f238d6398f396137e537e1379c363d3651358c33f2301d3140338d31cf2f;
// music[7192] = 256'h3e310c31742f672f042e822c372c532a4929d528b0281f2a7f29082915283924;
// music[7193] = 256'h762423273a266b25af248923742407244725e4255222a12def3feb4251426e40;
// music[7194] = 256'h643d0642d2457e43b33ed53c3d3c9539333a043797317233352d8f1bf214df16;
// music[7195] = 256'hdf12b81866211c11b800330096fcfaf8a4f68cf302f51af522f4cff5c3f581f4;
// music[7196] = 256'h53f4a4f4e9f593f54bf308f360f251f032ef33ee91ed59eb83e714e59ce49ee4;
// music[7197] = 256'h6de15edef1dcfcd876d7a2d758d462d34bd32ccfdacd84cd94c9baca37cb9cc9;
// music[7198] = 256'h4dd5f2e0bce059e0a8debddc36de62de42dd7fda93d8d1d88bd71cd76ed65fd5;
// music[7199] = 256'h51d47fc8c1b8b1b691b968b89db860b81cb71db940bb90ba3cbbabbc52bbbaba;
// music[7200] = 256'h55bb45bcacbd4abce9bbfdbb47ba72bc6ebd88bb1ebc9ebd4dc057c09abe11c0;
// music[7201] = 256'haec063c1d9c17fc1b1c32dc465c401c6f0c502c6a0c504c6e2c615c78dc908cb;
// music[7202] = 256'h8dcabbcad5cbcbcc7bd16fe1b9ec26ebadecf3ecf0ebedee46ee12efb5ef6aee;
// music[7203] = 256'h0af069ef10f00bef38eb2eeaeedf45d5ffd6fdd6b7d5c2d6c4d463d400d723d9;
// music[7204] = 256'h33daa9d995d967dbd5dc1cde59e080e0a9dfafe1eee2b1e116e3e8e421e36ae2;
// music[7205] = 256'h8be4fde557e58de5c5e72fe7b8e624e947e94ce929ea26ea7bea56e925e98dea;
// music[7206] = 256'he7e906ea06eb15eab5ea16eb46e97dedadf000f2ad009709a4050409e209f208;
// music[7207] = 256'h040d2b0cd10be00bc80ae00bba0bfd0b7a08b006d606b8f7baeb51ef4aeeb8eb;
// music[7208] = 256'hd7ecdaea6ceabfeb4bea10eac7eb8deb8aeb11ec08ec28ed93ec83ea17eb16ed;
// music[7209] = 256'h53edefeb1beca4ebadea3eede8ede1eca9edbaecdcec8aed3cec79ec11edfaec;
// music[7210] = 256'h70ec1eec1fed05ed3bedaeed5eedd8eee5ef40f068ef8bef1af35bf121f6b608;
// music[7211] = 256'hf30f8f0dff0c510c6311ac115310281b0f211021aa232523d72114204e21b21e;
// music[7212] = 256'h7d0dac023f050e068e046101c2ff77023b03c101a1002d005b0122022e012a02;
// music[7213] = 256'h1a043c036002f601c501a103bc030702dd01000266027e0213018bff32ff4801;
// music[7214] = 256'hef0271012f01e6012e03dc021cfbb4f987007600f202360762052d073509dd07;
// music[7215] = 256'ha808a1070d03190603118b155a197b1c68181d18e4149f0fd610830eb20e1f11;
// music[7216] = 256'hcc100613f01388190b1f411436021efd3e07600db80e6617671d6d1a1713950d;
// music[7217] = 256'h610b3c085c06fb03bbff74fd3ffbfef8e5f611f539f4f7f3daf424f56cf539f6;
// music[7218] = 256'h55f6eaf756f936fa1efd01ffb5ff4e027b04a605ae0757094e0b180ddf0dfe0f;
// music[7219] = 256'hca11d312e214ab16fe18451c7b1d191d41255534ba39eb39fe3ddf4003438f43;
// music[7220] = 256'h44432d4406441245624444423d420e42b9448740c731842cf32d322bce29a228;
// music[7221] = 256'h0c2851293c29c929272ae329c42980289828cb28802835299d2870288f28d127;
// music[7222] = 256'h7d287328d327f2278d279927e827a8279c27e9277727e8261a27ed260c27c526;
// music[7223] = 256'hb92581252b2569243b232723332309222c237a23a8222d225721f62a0a373737;
// music[7224] = 256'h99379f39b737fb37d938a9371e366235a13424322e310e312930ed309d29221b;
// music[7225] = 256'h8417551723127b125612f80e930fc90f9411ff132d11960fad0fde0d5c0d3c0d;
// music[7226] = 256'h140c7a0bf90ae00a7f0b9b0ae308ab08a00a500d4d0c9109fa087807be05c504;
// music[7227] = 256'h9b035203810207027e0246027d01ccff9e02fd09340ab8057a057e03bcfeb1fd;
// music[7228] = 256'hb8fa3ef98d05dd10f91002144f17ed15f71622184b177915fb137f12eb0e230e;
// music[7229] = 256'hf70c800afb0a14001df04bed70eaf7e4e4e4b6e2a6de7edcdeda86d98ad713d6;
// music[7230] = 256'he7d4e0d2bed1d6d06dcf6cce11cd76cb36caaec8e5c6b4c5f5c4e7c30fc342c2;
// music[7231] = 256'h0ec16fc0dabff0be55be9cbd4dbd9bbd56bdccbc9dbc16bce3bbc9bb28bb94bb;
// music[7232] = 256'h55bceebdf8be2ebdc9bdacbc10bdaecab6d4c4d4dad60fd8fdd88dd9b6da29dc;
// music[7233] = 256'h4fdaeee2c2ed38edaaee9cefb0f154f553eac5de69de2ade70dd77dd56dd35dd;
// music[7234] = 256'he4ddd6df67e0f4e02be2f8e241e4d0e4b0e4ebe43ee56ae5abe512e627e680e6;
// music[7235] = 256'h30e7c5e76ee8f4e8b4e96beaadea94ea71eac6eaabebbaec13ed38ed20ee0fef;
// music[7236] = 256'hc3ef47f0e9f081f10bf2c6f3b2f55af516f569f6e7f4b2f7b605cd0e760e3e0f;
// music[7237] = 256'hc20fbe1084129a1207132c128410a30fd40fbf10a70fff102b10430386f847f8;
// music[7238] = 256'ha0f837f902f9b1f7d5f7ecf5edf624f6e5ea0ee5e3e6d5e6a5e704e77fe63ae8;
// music[7239] = 256'h44e879e851e91dea92eaa0eadcea00ebb3ebd2eb27ecd5ec9cec78ed72ed20ed;
// music[7240] = 256'hd5edd1ed39eefcedabedc1ed2ded4aeddcec30ed3eee1dee84ed30ed29ee4fec;
// music[7241] = 256'h28f04300b506fc03b006e606ec061009e808a80921080506230617060207c005;
// music[7242] = 256'h1e075007f9f821eedaefe4eeb7ede1ed4feb66e9b8e809e995e9c6e92eea7cea;
// music[7243] = 256'hb9ea7eeab6ea88ea06ea9dea6fea24ea1beaade998e939e995e98be9a0e862e8;
// music[7244] = 256'hfde748e838e879e79ee768e7cce74ee8a5e8c3e9eee905eae5e9eaea0dee3def;
// music[7245] = 256'hbfefafef92ef36f0b1edfbf43006be099806df07ba060807eb08b90a3b0b6407;
// music[7246] = 256'h650640067b057506c904b706410220f172ebbeed50ec23ef99ef49e810e399e5;
// music[7247] = 256'h61e9afeb93efaaf1c4f2daf361f36ef3d2f130ef9fec85e99fe8afeca9f1e0ed;
// music[7248] = 256'h3ee9e1e8cae4bce327e4cde2dbe4e7e5f7e7cceae8ed52f572fa93f47be9e7ed;
// music[7249] = 256'h08f9fbfacf03fa0abc0a1d0e660cc10b390b4106230f341af817b014e612e610;
// music[7250] = 256'h0110fc0eda1179138b10d211c812f11289152216a3194814e70505051608cb08;
// music[7251] = 256'h750bea0b820e670e6f0c2e0f0c111d13921517172319771a5d1b5e1c021ea31f;
// music[7252] = 256'h29216922da22d7245126ef263028742802291d2a242b342cf02cd12dc22dab2d;
// music[7253] = 256'h462e8c2e4a2fe02fd72f30309e304b32a733d1329d32ee312c3147310232063d;
// music[7254] = 256'h5f49d04894470348bd46b54695456b47ab49e7484847814852531c598255e755;
// music[7255] = 256'h0c4d593e693d6b3f043eab3e203ead3de63cc438a5360a379d369c36cf36e436;
// music[7256] = 256'h7b36df354136223675353c35e8346b344534f3338133693372328c31fe302730;
// music[7257] = 256'h5a30ea2fc22f1930252ff12e422ee12c0f2c372bdd2afc2a872c7b2b3d29f52a;
// music[7258] = 256'hc92b6f2c292bc4296b34e33ddc3ba03a583aff38c838d838a139f4389a38053a;
// music[7259] = 256'hc73b873dad397b369c36e929791b111a091aa519a5193919d319f915ea10b20f;
// music[7260] = 256'hbe155c1bac0f6a01d7fd46fa63f8b2f79bf476f30ff3f5f2edf370f42bf594f5;
// music[7261] = 256'ha0f44ef47bf400f31ef263f11fef02ee78ecbcea53ea9de8c9e677e55ee3d0e1;
// music[7262] = 256'hf1e1a5e104df9bdd82dbfad895dadad77cd7cde4deeb0ce8d8e77ce7fbe56be5;
// music[7263] = 256'h15e398e1ccdffadebedfebdd6ddc38d98ad719d89acb1cbfdabf36bf26beefbe;
// music[7264] = 256'h45bf39c082bd4abb3dbaebb72cb80cb927baeeba5fba6bba53ba2cba9bba19bb;
// music[7265] = 256'hebba9cbb4fbd11bdbcbd8abe9fbd72bed6be23be79be78beadbe6dbf31bf59bf;
// music[7266] = 256'hbfc038c110c267c272c28ec51dc6f0c469c689c7dcc92acbe5ca11cc82cc74cd;
// music[7267] = 256'h76ce27cfd4cf45cfc6cf02d1c7d1cbd26fd453d6efd7c6d622d4c0df1cf215f5;
// music[7268] = 256'ha0f3dff508f619f6b1f5a6f6e3f75df6d8f5cef7a8f71cf68df762f88ef8bff9;
// music[7269] = 256'hdef912fbe3fb66fc73fb0dfc89fdc5ee2bdeccde94e075e1e3e495e580e431e2;
// music[7270] = 256'h53e131e366e402e480e721edf2edc9eccaebdcef42f6f4f4d9f39ff37ef230f4;
// music[7271] = 256'h39f00fed60f32ef961f9dff2ceebf7eccfeff4ef50f1b0f239f3b2f198f086f4;
// music[7272] = 256'h5bf7fff78df7faf26cf130f27df226f5cef4eff332f5cef3e6f155efaaee12f4;
// music[7273] = 256'h37f5a5eefded81f348f67bf6cbf490f26aef86ee60f493f618f5e2f69ef865fb;
// music[7274] = 256'h2cfb6ef698f3c7f5f601360fb61230153e19d4164a0f290cec0f301581164f12;
// music[7275] = 256'h2d0f2611bb154d19fc15a610710fb50cbb0cae14051cdd1dd41a7f13c805fef6;
// music[7276] = 256'h3cf48af9ea00f1073c0346fbeafa1efad1f929fb1dfbc4fb6bfbc1f870f7b1fb;
// music[7277] = 256'h27fab8ec95ea26f3cefac8079c07dafff505ef030900e009dd113b18821a2319;
// music[7278] = 256'h0d19c6144b13201018072603e00306074d05490246074e0407fa0bfb8d036007;
// music[7279] = 256'h1c069209d10dd909e60ac314c11bb81f491e431b8f20d0286e3122383f35892d;
// music[7280] = 256'h522a582c7e2f87357b3a5c3d4041853b7038d23a88357c44415c8260b8641665;
// music[7281] = 256'h5860c561d3620e65635c9d4c7953de6131617c613263a85dae5d1a62b161b35f;
// music[7282] = 256'h3f617d653161b7598d558948a13e964579490b3d7431ea2b67239f22b6289e30;
// music[7283] = 256'hd03d7442f93dd332b525fb27552ee32e1b30a02edd2d5730c134fc3901361d2d;
// music[7284] = 256'h0a2e8b2a18217d25952ae52b722c33238a22f1244f1c7315550e120fc5154914;
// music[7285] = 256'h7b18ef19c60ecf098b0878003ef778f3c5f51ef7abf5a0f57ff276eb34e783e7;
// music[7286] = 256'h0de9dfe539e0e6da69d6edda2be004db6ad9a9dfbcdedad89ed63dcda7c44acb;
// music[7287] = 256'ha8cb13c699d239e58aeb1becdceab9e375ddced927d5d4d7ffe1e1ec03f1c0e8;
// music[7288] = 256'hb3dc49d6a9d80cdcead9ecdb67dff5df31e32de3f8dea0d95ece1ac8bfcda4cd;
// music[7289] = 256'hc1c50ac661ccd1cb14c8f6ca7bc905c59dc64fc0aebd21c8bece33d561d6dcd3;
// music[7290] = 256'h15d691d019d1eed695d213d5e7d6a8cf46cb2fc5d0c44dcd98d348db93df0cdd;
// music[7291] = 256'h05dc6cd7bdcf9fce42d65ee077de98d889dc1ad93ed19fd544daa8e039e6bdd7;
// music[7292] = 256'h72d004dc19dbc0dc75e79de235dffae619ea5ce41ade48e146e634eaa8edbbed;
// music[7293] = 256'hd8f259f540f4bdf33ce8f0deffdfc9e181ec16f53cec4dee3a011b058205670d;
// music[7294] = 256'h6c10f01a3821251b9e1c8b195e11120f1a096b06980bfd0e14136f183d1bf119;
// music[7295] = 256'h910cd800cf057605bcffde0216074f0afa061602c5047b09aa135c1d071b2712;
// music[7296] = 256'hc40d8e10d1158e1f99256323bf24812a112c6026af276f32103637363f36cb33;
// music[7297] = 256'h7330813142385b37c9329734b339053e8a392b35143580364c41024300323529;
// music[7298] = 256'hce2f733b2e403d35dc328e3f7a3fec3b7d3c793b413b9035233bc53b952a8037;
// music[7299] = 256'hb049c4408140a24b4751634910408042893faa3dd3424e3bdb379641ce3f0942;
// music[7300] = 256'h6f53755c985c5552fc48cf4e9755805bea5493477d4a0e4a0f48b04ca4460e3e;
// music[7301] = 256'hdf407741d43b8140103d752c0d2b342c142e942cff1759098203da00bc054b03;
// music[7302] = 256'h4d018b01ccf958fa34fdb4ef55edf1f7c2f1d3ee27f708f708efbbe3b7e393e6;
// music[7303] = 256'hf9e124e987ebbadd48db11e177dc52d7c4da99dfe0dfc5da94daaaddebd985d8;
// music[7304] = 256'h3ed497d312e14ddd16cd9ac823c3b7c0e9c505c877c630c336c7dacc23c3ccbc;
// music[7305] = 256'h16c471c72fcb18d0f4cab5c0c7b9d7bb26c2ebc626cb4fca5dc96ccb69cbc2cc;
// music[7306] = 256'h58c74abc6ac001cbbdcac9c98dd50de8aeeb34e114de4ee3ede596e344e3c9e5;
// music[7307] = 256'h9ae80ceed6ee00ee15f055f2b6f478ed8cea0ef2eef398f823f235e410ee10fb;
// music[7308] = 256'h72f4e9e3d4dc65df3dd8ebd486df11e56be367e483e3d8de3ad8c4ccaacb7cda;
// music[7309] = 256'h60e77eef2bf12febb2e5e8e94bf083ea05e619e81fe604e329df57d610d00cdb;
// music[7310] = 256'hefe4a8e60eef06ef77f5e9006bf31ded04f624f474eeffeed2f0ffee5ff082ee;
// music[7311] = 256'hc7eb06ef90ea64e99fef14ed79e87bee8ef6d7f085f027fb3e00b6074a0a2e03;
// music[7312] = 256'hfc0215086b0a3e0cba10f112da11bd0f9c183e22c4163314cb1ad81e12392946;
// music[7313] = 256'hfc40c7492a4664396439b13d4946984bcb4b48546355ac490f49be48154bb958;
// music[7314] = 256'hb754884eff52594ea14d69539d55a04fe143ce3f3d3c2e344f31da33c1331330;
// music[7315] = 256'h5b304c330336db335d2bd52a3633a83537323c37303c6c352e2d562578279232;
// music[7316] = 256'hea3529394333f728b72c472b8d2c2835e130382e3f2d0128a824101cce1d2b24;
// music[7317] = 256'hd716d50f6b111509600b8e12060b980188fc05fa02fb6ffbc8fa51f768ed82e7;
// music[7318] = 256'he5ea3bea89e394dfbddf37de57d851d56ad181d1f4dcc8dd8ed96ddbaad7e4d8;
// music[7319] = 256'h03d6dbcd4bd341d38cd995ed3eeaffe1fae8eee81ee47de2abe590edbbed69e5;
// music[7320] = 256'h60dea3dd6ce222e5dee637e6e3e20ee890e6b7e134f0abf249ea75f213f0f6e1;
// music[7321] = 256'h79dc96ded7e115db26d5c7d800de06dfafd6f1d25bda65e2d0e6ece6d0e436dc;
// music[7322] = 256'hacd366d3a3d07ad3bfe048e70be6ece156d807d450db3bdf16de0fdfafde0fe3;
// music[7323] = 256'hfee922e663e051e5d9e52ddd1edd80dfa2dd7adffae116e5f0e480e210e33fe0;
// music[7324] = 256'h47dc53dc50e1c1e3d8e440eed8f107efc8e8a8df1fe4b6e606e681ed50ef34f2;
// music[7325] = 256'ha7efc7e42ae94df1aef364f884f613eedff3ca0279fe02feb011bb0cba01310e;
// music[7326] = 256'h17024deed0f7fdf732f4cbfeaf05c40b510de60a250d3d0de40d3f0de00a040c;
// music[7327] = 256'he20c520ba908fb0a1d0846f7a2efdcef4fec7df46ffac0f4a9fce7ffcdf87200;
// music[7328] = 256'heaffb0fe180c4c091906f40bcc0bea125b1771127f115d15bd1dee22d41ffb1d;
// music[7329] = 256'h4f22ca20aa177217451b861dab23362940307d339e2ac8239e2632289e25e228;
// music[7330] = 256'h533065357d34af2a6f2c6b370b302e294c30d835153bc53c2334cd266023652b;
// music[7331] = 256'ha22ddd2e5a353537ff344430c02ecc2d0a27052d6d37502ccd23512d49317b31;
// music[7332] = 256'h3c30c923d82adc477f4997388136773acc410f4a7a4d804d2e42013d0e438b3d;
// music[7333] = 256'hbc3d8e429a3b49396f374a353b34df2dc22e42291e20df22ff104df746fa1401;
// music[7334] = 256'hcafc25f725f282f275f1b1ec13e957dd50d853e495e61ce66eec98e3b2d5d9d1;
// music[7335] = 256'h0ad43dd776d07cca8acafbc1e8c214d0b3d078d1dbd37cc85dc4f3c8d7c4b5c3;
// music[7336] = 256'h0dc8e4c9aac61ebf97c05dc38ec092c5d4c526c28cc409c235c539c82fc0babd;
// music[7337] = 256'hdcba9dbb4cc6bdc30dbe7ac7e3c93dbd77b758bec5c9fbcf85c7a9bf42c252c3;
// music[7338] = 256'h73c22ac612cb1fc928c8edcad3c69ac3d0c427d2f3e4fce12be01fe6e5dd25e1;
// music[7339] = 256'h18eb72e3e3defadfbce1beecdeed43ea4cefa2e8dee276e51de80ff1fded54ec;
// music[7340] = 256'h2af32deee9ea14dcf0cb22d2ded4a8da9fdc91cf4ecf73d677dd48e382e33ae7;
// music[7341] = 256'h9ee80be6aae2abdafdd6e0d57dd322dcdce53ce78eee63f3e2f3d6f2fee136db;
// music[7342] = 256'h04e6f9e7d4ecd0eb5bdf9ee5c3ed81ec96f948041804df074805a2048d0c3c08;
// music[7343] = 256'h87015cfd6af563f9b2fb9df8ba029206e9079d09cff956f8fdfe7bf8a9009b08;
// music[7344] = 256'ha60695042e05d0141e183a11e617c719b81d5621f41d39213625fc2847294a27;
// music[7345] = 256'h52313241984dba53f450844759449a464b46064da5538555af59f1583959e35a;
// music[7346] = 256'haf559a50b6546f62126933642960cf57a1508254054fc8418e42db466c4a974c;
// music[7347] = 256'hc243863f73430943e642224524426d3e4d4339439d38db2cb928eb346937d32c;
// music[7348] = 256'ha1314f340c29ff204d206a22be248a25092736300a32512fc930951f8812c11a;
// music[7349] = 256'hff1db920db214b1da41b0819cd114d0ca60ce3092309f80a230503067703d7f7;
// music[7350] = 256'h4bf70ff5c3ef77f2c4f0f1eb05eb3eeb9cea44e59ddecfdfe7e2f4dd23d8efda;
// music[7351] = 256'h27de6ed836cd4bc550c7e3c9cdca00da1eedb9f1d5e701de88e2c2e654e39edf;
// music[7352] = 256'hf8dbd1ddb3dfbee0c0e0fad607d350df14e80ce345e055e081db8bda25d833d8;
// music[7353] = 256'h35d633c5d7c43dcdd5c0cbb91bc240c6cdbf1bbeb6c882cc75c814c77ec51ec3;
// music[7354] = 256'h23c3d1c5cfc9b7c8c9c47cc87fc96cc87dcc4ac394bea5c84cc8bdc97bcdfbc9;
// music[7355] = 256'h57cfc7ce7cbf10bf15cde2d0f8d067cf23c7c4cae8d0cccbe7c801c7d4c998d2;
// music[7356] = 256'ha4d431d275d26ad419cfa8cd0bd610d3a2d168d877d231ccc0cf12d44cd564d9;
// music[7357] = 256'hdee00bdf53de0ae01adba9e0b8dfdbd0ced456db3ada5ae30ae150dceff4c408;
// music[7358] = 256'h8d062b053cff8ffc7d032f0296f96ae9dae08aecd4f3b8f85b03870ce0167117;
// music[7359] = 256'hb010320bf907e612cd18ff121d18b30f80f459e7b7e307e540ec76ef98f62b02;
// music[7360] = 256'hcc078d06bd0123fe48fffa05b6051200bb07b30ea10d98102c0e3c0a88111916;
// music[7361] = 256'heb118716121fac204e28462be4223d20b51ed420b5227b1f862500250523982e;
// music[7362] = 256'h9c2d2f260324ef233d2d8430722fba31652cbb2cb72ee02b6f332b37c2331d33;
// music[7363] = 256'h3c30de314931d22bae2cda294d28ec2f75308e2f2539223ac92dbb2a912e3a35;
// music[7364] = 256'hd2420c4540416042393fcc4669559f556654c656c352084fe54e4850ed548355;
// music[7365] = 256'h4b539e55a953be4d584b4e4d4a536b524549eb45ec4bbb4d6a45c041d2398e1f;
// music[7366] = 256'h6411bf17dd152f0d820a1d0ce60f9e104810340beafd4ffd8602e3f959f170f0;
// music[7367] = 256'h3ff4d6f3e3ee48ef91eb4ce79be47dded4e3a0e75be246e6b0e9b8e66fe327d9;
// music[7368] = 256'h35cdfac755c7e4cea4d378cd94d491dd7ed4c9d1f5d3ecd2f2d2cecbb2c94ecc;
// music[7369] = 256'h62cb67d0edcff8c98bca2fcacfc5e4bc0fb728b975b8f9ba61c17bbffabc80c1;
// music[7370] = 256'hd3c54ac1d6bb3fc294c898c4fdc1a3c2bdbcd2bb86c50cc87fd080e2f4e5a1e4;
// music[7371] = 256'h18e04dd784dcffe3c8e49ee999ec69e54ce494eb88e709e724ec2ceb6fed07e9;
// music[7372] = 256'h80e5c3e5e4e0adebe6f276e58fd670cca2cd77d531da45dd75dffadc30d8dfdb;
// music[7373] = 256'h8adb86d74ed809d390d367df7de71ee4b4db27d521cec2d3b6daafda8ae2e2df;
// music[7374] = 256'hdddd51e860eca9ef64ec0de3eddd01ddf0df27d528c7b1cc4fd59fd4addbeee7;
// music[7375] = 256'ha5e753e905ec8be842efc4f122ed89eb07ea4cec67e98de47feb41f467ee81e2;
// music[7376] = 256'hf1e4dae83fec0ff4c2f594f951fae8f981fd27fcb303d709dc0a8b10cd080005;
// music[7377] = 256'h590d2a0d581247258e34123b574251423b3aad3bb23bfd3aab41a63ed73aa743;
// music[7378] = 256'h464d584e634994474449244c674a3c477e4def4921466d55bc4d7a36af32ec2d;
// music[7379] = 256'h972f5637d332b8398843b53e5b3b2c35c52d50332d3a31359a2faf3382351a30;
// music[7380] = 256'hff2b412b052fba363639213529341733752cd1264121b41cfb1e4d2327252f29;
// music[7381] = 256'h022af520e72111294f229c215625e821a7225c1c6d15c6193b1aef19e818e910;
// music[7382] = 256'h940d690e5c0ba8064a03970295ffb7f70ff632f634ee80eafaeaece624e6fae5;
// music[7383] = 256'h07e247e474e528de45def6dcc7d8fde081db10d9e4f292f54be5fce5daeab9ef;
// music[7384] = 256'h1af036ee6bec7ce383e20fe6c2e5e9e70be330defae250e603e67ae24ddf68e4;
// music[7385] = 256'h3fe469dcece19edfa4c98dc953d089c721cfccd658d00cd4acd99fdb66d9c7d4;
// music[7386] = 256'h21dab2d997d5d4db4eda8cd4a2d449d121d0a1d546da81da81d98ed9c6d8d3d6;
// music[7387] = 256'hb3d019d049dc1edcbcd054d283d63cd4fbd07cd4a5e02ae3bfdd2adca9da8cdd;
// music[7388] = 256'h22e015e154e60ee583e548ebb0e45fdce1db89df9de6a2e7f2eaf9efa6e908e9;
// music[7389] = 256'h4dea95e5b3e935eae0e755ef19f6abf65ff04aec9aeee9ef1bf36df1b2e96cea;
// music[7390] = 256'h17f86508110bf2032605d00fc816e5158a12b90aff07701380144102fcfbd001;
// music[7391] = 256'h1bf9bff23dfc7202ab05220efd12bf0aa60cc219a40620eec6f144f737f96bf4;
// music[7392] = 256'h41ee1bef2deab8eccff35df0aaf197f802fb95faa0f70af598f639fb31044c0a;
// music[7393] = 256'h76055d059a0d1c12d9119111a618761d8614320d97117818411e7124ae20eb1a;
// music[7394] = 256'h22227f2a322ac225a128712c4827b42aaf328a315c2e8433e036ff270f268535;
// music[7395] = 256'hb833402c86296f28be277a2ae835bf34012b3b2b732d9b2e3e2bc727ef2ff836;
// music[7396] = 256'h81323a2f352a8122c227af25832063338647364ffe4afb3e593dc142f442d33b;
// music[7397] = 256'h963d9b41273d9a438149944856473a413e412a3f7b3f9943cd3fc4416f3a9b30;
// music[7398] = 256'h5837512d181a0d141d0ce106e20b510beb05c105d801730031020bfc7cf9f4f6;
// music[7399] = 256'h2af4d8f46fea89e2fde6c4eae1e7bce2e5e009de9cdc80d766cff8d4e3d520cd;
// music[7400] = 256'hb8cba0cb89caacc883cab2cca1c505c42dc5dfc370c6dbbf65bbb1c1f9c016c1;
// music[7401] = 256'h98c25dc070c2b0c0bcc1b5c4b0bb9bbb7dc012be21c2adbda0b637c164c625c1;
// music[7402] = 256'he3c0b6c055bf5ec222c1adbce6c2d5c626c4bcc38fbe61c236cb4ac57cc830d8;
// music[7403] = 256'hc1df4adfebd9bddcd8e509e4ebe2bfe54de345e6d4e815e376e518eb3fead7e9;
// music[7404] = 256'h99e741e81fea38e50ee879ed68ebe3ea9cdf3dd15ed6b0d956d51ed96cd754d3;
// music[7405] = 256'h26dad0da21d809df34dd6fd28dd0cfd36dd73bdb62dc81de02e380e436e380e2;
// music[7406] = 256'h46de79d740d698d968dfe6e44ee25ae0a9e8bdec18ebc6ef2fefdbe5f5e2bce4;
// music[7407] = 256'ha9dfd5d07bccbcdd95eb15f35ffc17fe26006e0335024002a6018004ac071103;
// music[7408] = 256'h7bfe3bfb24fc75fdacf58df3d2f99efe24031104f204470526014204810aea0c;
// music[7409] = 256'h45133d176817de175713671da438963dad34253ab9407f451c48d844e548354f;
// music[7410] = 256'h674fe84c4b4cfe5084529455de5c1b5946561e5e625f2e57ed537b5da460c54e;
// music[7411] = 256'h2b44ef481e4757464c48c947874ed54b39405e441e4b4445153c563a873d6a3d;
// music[7412] = 256'h573d59410649d748723edc3b4c3a6c3497389f3d5239e435f730b325df248b29;
// music[7413] = 256'h5922b81f1726ce2950284221d91d75226727d523221f1e21831df31d0f226b1b;
// music[7414] = 256'h411a5919b4121d100f0a4409e509ee03ff081d0b69008efd22fce0f619fbc6fd;
// music[7415] = 256'hb9f6dbf4b7f30bed2fec46eb21e889e7bfdf08dcdcdff9dcdde333f1f8ef9eec;
// music[7416] = 256'h64edb6ecfae96fe9e8eb0be65fe2a9ea18ee47ec28e7f4dcc0dc0be26edf3ce1;
// music[7417] = 256'h3fe5c6e09ee07fe2c8e05fe098d3bfc259c262c5bcc4c0c2a5c012c7c9c724bf;
// music[7418] = 256'hcac331c89ec38dc39dbee6bbc9c13ac31cc4f9c4dec6c1c8c1c312be5cc097ca;
// music[7419] = 256'h52c8b0bd91c26ac5a8c26cc374c40cc938c95bc648c4cdc438cba5c8cfc52dc9;
// music[7420] = 256'hbdc732c90fcb95c87bc660c686ca64cd2fca91c83dcf4dd113cc37cc0eceabd0;
// music[7421] = 256'h6dd2d9cf8acc59ce27da86dd22d94edaf5d2f6cf6bd68cd555d804de6dda49d6;
// music[7422] = 256'h0ed883da24e25eed3becb9ea84f3defcd50288003dfd89027b064a03ce023103;
// music[7423] = 256'hd6faadfd67085d0178f5daef3bf50a05c50c610b930b4417bb1b7a062af884f9;
// music[7424] = 256'h4ef7cef7e5f850f58af500f594ef82ee97ef35efeaedc0ead0ee77f493f5fef8;
// music[7425] = 256'h35f8d1fada01d6fc16fd6e07f50673031507a80c4810440fce108f13e911d415;
// music[7426] = 256'h9417b5147a19c41bf61e37216b18b7178d1b431df42584267f1fdc1f9127c42e;
// music[7427] = 256'he42d032cc62dd72ed92fe12fc62ef72e9d304530bf2da12e20376841f9402439;
// music[7428] = 256'h5f3418369137b02e672c1d352138e73b1139fa35f746184e8b4645502461c862;
// music[7429] = 256'h445ac358975a6753e551a35b1e5af45164555c5a665cf75c055ab15aac5a525a;
// music[7430] = 256'h5359c3556f5a3852df3907314030c92ada2551218d1cc61da122ef1da71a8e16;
// music[7431] = 256'h790b980d7d126d0fb109fc025205db01ecf6f3f668f88bf572f7b7f909f64ef4;
// music[7432] = 256'hb0ee45e334e47be515e0d1dd40deefe3e4e752e72fe192d92bdb1ad81dd453d9;
// music[7433] = 256'h6ddb25d995d73ed881d37acb98c93bcacdcd39d1c3d205d1a0cb72cfdcd419d2;
// music[7434] = 256'he1cfa0ce02cb4bcb56cca6c487c1ddc476c416c595bf8fbdd1c46bc582c48dc2;
// music[7435] = 256'hadc245cf3dda80dac3da11dfe0de34e1dde4b9de72da7bde8ee5aae455df2be2;
// music[7436] = 256'ha1e02be2ede712e74feb90ec1eed9cef4bedd5f0ffe6efd428d5ffd619d7e5d6;
// music[7437] = 256'h35d182d16fd53cd726dcc5dcdad3a6d063d62ed80bd6fed555d904d95fd2dacd;
// music[7438] = 256'h5ad243dc84de08dd87dd70dc20e0b9db9dd564dfebdc21d6b1dd85dc9cdda4e7;
// music[7439] = 256'h59e8a9e2a7dccfdd76e032dea6dc6cce1ac3eece52d50ad7f8df3de151e503ef;
// music[7440] = 256'h9fed2aeb0bf268f5a0f111edd8e7ecebeff2dde82ce39cec5df061f2def4f7f0;
// music[7441] = 256'h01f072f5f2f898f823fd9302fcfc52fc490e5a202328d02a82266921b825442b;
// music[7442] = 256'hac2c6431e2381d3dfb3a5b380c3d4040913ebc3f3141e5413147864f854f2c4a;
// music[7443] = 256'h754cc748b33abd2f142ce8321f369a35c23d383a562e81314c39233736331f34;
// music[7444] = 256'h14317a311335462fe52fa833692d582bf62d5d32163964390836c133be2c092a;
// music[7445] = 256'h1e31fd30bb2e6831d82d842cd62bbb2559254d28f828892b3d2ccb25bd26e52c;
// music[7446] = 256'h4c27cf281e2da1245e20a51ed91d401d68182a196d19df181319a1149a130313;
// music[7447] = 256'h3c0e2807b3febff9a9f88bf8f5f6acf38ff340fad5f905efb8eb49e659e7e8fa;
// music[7448] = 256'hf50172fe5bf985f1fdf4cef509f38ff57df207eef1edafefedee80e8cfe4ebe8;
// music[7449] = 256'hdcea6ae868edc3f242f2b3efc9ec30ee03e293cc59c80ac998cbc9d1eacf68cc;
// music[7450] = 256'h72cd97cf79cbb9c7a2cd5cd2a8cc92c4b5cc7adaf7d9ecd6d8d559d5b2d534d9;
// music[7451] = 256'h24df48da8bd729ddcdddeddb65d530d5efdad0d721d882da28d9bdd8feda5ae0;
// music[7452] = 256'hebda30d662dc8ad91cd78cda94d9ead862d75ed843dbbcd9e7d9dedc19df16da;
// music[7453] = 256'h88d78ce3eae59edf1ce2e8e11de62ae956e477ed15f192e94eebdae6cde527ed;
// music[7454] = 256'hacea56ecaaefdbec24ed84ef4afec40fd80e29092c0365fd3002dc053c070b0e;
// music[7455] = 256'h8c0c5606d10bca14d814fb107414d819c31753131606b0f699feb40c410c4402;
// music[7456] = 256'hf1f290f4ecfe12f737f5ecfadbf6c2f5c1f3b5f02beeece835ee02ed92e2c8e7;
// music[7457] = 256'hd3ebbce9b6eb12e96dec76f610f7eff68bfd05009cfe71ff87fe6902bc0b710d;
// music[7458] = 256'hc50c640bf907d40b0f0f7b0e6d1263170e1abd197718a01cc025b029bd25be23;
// music[7459] = 256'h3c23ba22f7244f24a0241a26cc24362a7b306d32913683333c2ea3303930b22f;
// music[7460] = 256'hef2fca2e7934ac367f38e63c66346e329635b62a5225f9263832fe472b4f954a;
// music[7461] = 256'h654553434c4258434e4ec14b23414845334624434f3f6d3b013e08400d43a446;
// music[7462] = 256'h0b4a574a0448204cbc4a7e485a41fe2f932eca29fa1fa226bf238d1fe9211e1a;
// music[7463] = 256'h8a18eb1c1f163a0e240edb074cfecbfd51fd76fdb1fc81f91bfb35f4d4ea3dec;
// music[7464] = 256'h18eb99e632e42ce07cdae0d899dd12df70dae6d43ecff5cc8dd0eed364d44bd3;
// music[7465] = 256'h7cce58c9dfc5c5bf18bf32c5b5c5c0c5c6c87cc837c814c317bd72be92bd66c0;
// music[7466] = 256'h26c47dbe83bf8bc630c9e9c8b6c8b4c7e1c259c13fc241c47ec7f2c875cef9c8;
// music[7467] = 256'h12c25cc6cbc04bc8c0de26e3c6de31deefe2a8e387e095e082e1dde64de313de;
// music[7468] = 256'he4e4cde63ae7bde887e8a3e925ea39ecb9ebc2eb21edb2f22af5bfdee2cd0dd5;
// music[7469] = 256'hf6d5b1d175d327d5e4d255d508d8a8d3bcd751dea1da02d849da7eda71d707d8;
// music[7470] = 256'h62d664d229d687db86db95d6aed676dcabdc60dca5da50dd8fe631e187da6fe2;
// music[7471] = 256'h89e26ddd94e446e85de57fecbff190edbee854e567e442e253e52fe6d3d596d1;
// music[7472] = 256'h4ddf53e40ceae8f5eefc9400a1032906d905ac05ae060b02d80027054201e1fa;
// music[7473] = 256'h6af773f788ffaf009efa0c020e0a0905cb025a076316482b5f2be925e72cd22c;
// music[7474] = 256'hc22e153756352532fd35ff3da0400c3f2a447d455a45c34c29533c593659f656;
// music[7475] = 256'he45ba557b1534856bc4b07420841fb43074bc84713440848af49d34d564c8d44;
// music[7476] = 256'h7c45af486e4542420243f53e833ddc46b7474f41f9418842d23e8538c936893e;
// music[7477] = 256'hdc40f03c3c41dd408938ae35a834703d6846333bec30c22a4823f422ad202a22;
// music[7478] = 256'h0526c9201a23c4282d23961ef11ff920501f4a21b928ab21ad16eb1ae8183a17;
// music[7479] = 256'he918f40fbf133115130a0d0b760a8d0a800ac5ff51fc45fab1f723f7ebf199f1;
// music[7480] = 256'h4bf036f25eff1805a7031c02dbfacbf362f4f8f5e7f28bf325f931f723ef95ee;
// music[7481] = 256'h4df282f3c1f158ebe2e7f6e7a3e9b6ed97e8bde468e5ced712cacbc7d8c728c6;
// music[7482] = 256'h91c494ca75cc86c5c8c26fc1e7c344c3f1b947bd0ac53ec32bc1b1be2dc0c6c2;
// music[7483] = 256'h63c0fcbea2bc40bd4fc084bfecbba0b746c0d9cb21c728c2bac1afc08abfecbc;
// music[7484] = 256'h21c27ccb2bcbb9c5bac2a7c07cc212c7d1c43ec6f5cc88cb6fca79ca94c876ca;
// music[7485] = 256'h8ccd2ccfb3cbfdca8fcecccc18d01ed4bcd2e0d5a9d4ded06cd548d77ed18cd1;
// music[7486] = 256'hccd8b2d64bd35adbf5ddaddb97db22d744e3affb10fbc1f391f84ff8c6fc6100;
// music[7487] = 256'h2af413eeb7f476fcaafe9ffe7f0211ff7bfcab04bb08160abe07f2000e017103;
// music[7488] = 256'h930110f481e0bfdc88e17ae6ecf190f95ffa7ffc54003504f10077f916f840f5;
// music[7489] = 256'h11f1c4f3e6f44df14cf110f643f40cee90ef72ee0cf085f9e9f573f29ef686f7;
// music[7490] = 256'ha8fd93fec2fd5004be04af07420bcc0afa10a1122210b311c0136a17f11ab61c;
// music[7491] = 256'hd41936173920e928af256a222124b425c82b3e2fd229132b962f082f0f2d422e;
// music[7492] = 256'heb3577333730ed3ae13a04365737f935783461334439c53ccc37d839eb3b5342;
// music[7493] = 256'h4d4ed84e844f2c533152c952714f3a4c644c7a47224eb45914542e576a5f1f57;
// music[7494] = 256'hfe5443570a541556435a795a9657125cfb5be74ae34303461e448644723fbc3a;
// music[7495] = 256'h9c3a7a34e82f4b2f862d002da62cfa282a21fd199716a4158d15090f4007a00a;
// music[7496] = 256'hcc0dc008b8038cff2ffe08ff65f94ef431f91cfafef4ebf7b3f5b7e908e91eec;
// music[7497] = 256'h7ce5a2e21ee637e354dda8def8e2e5e0cfdc75debadd0ad949d6e7d254d31ed5;
// music[7498] = 256'h2cd65dd652cdb0cab6d187d295d45bd637d2e9cc89cbf0ceb2d039d2c4d046c9;
// music[7499] = 256'hd8c8d3d1fed57bd04fc8f4be6cc73fde4bdee4d7f4d9d9d8afdce2da03d7e3d9;
// music[7500] = 256'h7fd968dbb2dc7edcefdef5df10e1c7e08ee28ee270df05e433e41fe016e71ae5;
// music[7501] = 256'h1dd430ce94ccf7c9d0d295d229ce7ed768d6a7d1abd4ffd096d442dbead518d6;
// music[7502] = 256'h63d82cd6ecd849d938d894d51dd274d8c7d7a0d178d3ced19bd113d3e6d2e5d7;
// music[7503] = 256'h76da3bdbf7df70e264da2ad32ed76fdca9e2c2e287dd1fe3f1e6bbe6a6e9e3e9;
// music[7504] = 256'h20e76ee49be58ee13bd399ca68d288dd2bdc38e002ec95f1e6f7cbf6eef0ddf0;
// music[7505] = 256'h6cedeaecc1effeec78ec4ff118f2fbf0b8f123ef1cf26af50bf4bf02ef111313;
// music[7506] = 256'hcb174b1ae716cd165d1ad01f86211c211b240b26bc2a7c33f933cb3204356035;
// music[7507] = 256'h423a0437f630623a543f114282413f2e2126b92d1031fc310030043010321133;
// music[7508] = 256'hee3457365d39ed370734a831862e73332635d131bf34272f5e2e313a7535fe2c;
// music[7509] = 256'he4312331052e0e312c2cd5294a34b234a32f70330a31ab28b526492d5d344232;
// music[7510] = 256'h012f312e5c29d226fb28532a7e298825c223af27d528f127c12c3e31f42cec24;
// music[7511] = 256'h562133234b28bc28ce252525b01fba1c191c8915b7155d13e90c0a0f6a0d9009;
// music[7512] = 256'h9805ae009dfe9afb43068a113909d105280a3c096306b20003fbcaf8e0f7f1f6;
// music[7513] = 256'hcaf650f647f50bf6ecf54af134ecaaea5be93ae756e6b9e6d2e804e658dcabd3;
// music[7514] = 256'h76d282d3cfcd8ccefad392d23dd564d48cd1ffcf86c670c964cf99ca27cd88cf;
// music[7515] = 256'h0bcf35cde0c69fc79eccd7cc45c628c5c6cf1ad639d9c6da43d6a4d4aad25ccf;
// music[7516] = 256'h51d2bed756d993d686d656da0ad874d12bd23fd973dae9d880de83ded5d78fd9;
// music[7517] = 256'h24dc14dd6cdf8bdf3be023dd6fddcbe348e2f1e1ebe16ade04e166e2e9e2f5e5;
// music[7518] = 256'he1e7ace848e755e57de181e392e991e72ce770e6a0e86bf93f0379036a094208;
// music[7519] = 256'ha50194040a061504e508d50db30fc00866008906350b440a6e0bab0be20d6f12;
// music[7520] = 256'hfa1a5016230af910fb0a3af6f4f32aee66dd7add69ed36f34ff76e0390fd34f7;
// music[7521] = 256'hbbfbaaf378f2bff778f426f46aefe5e8c8e682e59eea13ee82ee2eef81ebceeb;
// music[7522] = 256'h74f053f3c1f6befc66ffbff931f7edf8d7fb1302ae012a014a08e10f78143a12;
// music[7523] = 256'h4b14a71bd51b3f191919991eaf20d81e04261126152070263f2d3c2a1624fa24;
// music[7524] = 256'hb12819287c2bfd2e192b3b2a05309d30802aba28bf2b8c2fd831c230d42d3028;
// music[7525] = 256'hc02875383648c64dee4fcf4dda45754009447c4d0950104b2848354617491a4a;
// music[7526] = 256'hf1442e4dce518b49764af145c53ec53f213cde409845dd385e2e4d2d772d7e2b;
// music[7527] = 256'hba2c762ff22a1d29842a33296f295e27dd23ad1ee918d7189d185917fe139c0c;
// music[7528] = 256'hdc09760749018d006904eb0104f8fff2bef478f445f335f302f2f4efc9eab8e2;
// music[7529] = 256'hfee0b3e4f6dfc1d72dda5ddd30da41da9cd73ecf7dcd13cf0fcf90cfe3cd1ecc;
// music[7530] = 256'h79cbafcca8cc70c861c958c837c08cbfcdc2b1c3c4c564ca49cb9dc3bfc16ec3;
// music[7531] = 256'h9ec30bc812c4a9c098c348c4a5ca8ec823c91adc2ee1c1dcb0dff7df39dd49db;
// music[7532] = 256'h2de04fe344de82db76db23e0a5e3eaded5df7ee6b0e55be2fde217e5e7e9f7e7;
// music[7533] = 256'he2e01be67ae0a1cc9dcba6ce53cbbcd1acd899d755d3c3d1aed420d666d056ce;
// music[7534] = 256'h9ad749d840d41ad851d33acf50d3cbd4ded9a7db26dbe3dd18da67d900db8dda;
// music[7535] = 256'h57dea9d981d469da18dc79da33ddccdeccdce7df95e330dcebdbfce239e04be3;
// music[7536] = 256'h99e7b2e1fde710f590f2eaea1ee823e7b5e878e970e3e9d8dfd525dd57e183e4;
// music[7537] = 256'hc8eb0bf1b3fabb05e807cb08030b33089200a4ffad0419ff87fc5f045000ff01;
// music[7538] = 256'h3c14d91a801b181e881d2b21a32209252c29b627132b012b1429f53194346432;
// music[7539] = 256'h90351a38583b613ea53f85435d4823499c4899429738d839173ac236a33e0341;
// music[7540] = 256'h1c3e2642774364425e45da482647a4431b429742ce463746074303441344ec46;
// music[7541] = 256'h74474c41cc3ebd3fd84393464e4442440941693d9d3d3b3a7e3d4841173ccf3b;
// music[7542] = 256'h833a4739bd3b7b379d3b7941033b623b9638f22a83273f27a223d324af246d23;
// music[7543] = 256'ha7250a261a236b221c28b627b020ad214f20471dc61e391a2c19e919be152515;
// music[7544] = 256'ha613b50e59093a09b90728ff9d07fe16a1147310d00f840b420910092b051302;
// music[7545] = 256'h7600fefa4df972f9b0f6ecf723f873f37beecdec59ec7aec14f03eec98e711ea;
// music[7546] = 256'h5ddc6ccb34cc51cdd6cd7fcfa3cd44cd14cbfac809c7cac3efc507c8f7c69bc2;
// music[7547] = 256'h77becec155c2cdbfa6c102c4b2c392c09fc28fc4d7c04fc012c063c019c06dc0;
// music[7548] = 256'h9ec34fbf45be27c382c0a9bebec0fbc293c213c136c473c56ec4ccc5f1c53bc7;
// music[7549] = 256'h99c881c571c402c81acab6c96ac7afc687c64dc53ac84bcb3dcd9dce06cc7ecb;
// music[7550] = 256'h83cd64d1cad38cd334d3afcfcad158d5f6d269d590d67ed3ded310e02eef07f0;
// music[7551] = 256'hb3efccf0bfed3befa8f339f4deef47f51cf94af2c7f5b9f788f9f0fd06f69ef4;
// music[7552] = 256'h0cf9f5fa180076029d00d6001309b1ffade616e467e6a9e1ebe577e670d94ad1;
// music[7553] = 256'h96db79e2b0e5b7f15ef684f8bdf9aff395f552f8d2f391f0a4ee7cef66f240f3;
// music[7554] = 256'hcbf1feee1ff08bf1e3ee66f294f8fcf656f589f8b6fcd5fc64faadfb43fe5e00;
// music[7555] = 256'h3f055e094b08c40a47127c12bf1219171d19cd1ac9193c1cc91f131eb8210223;
// music[7556] = 256'h821fa221732651293c27ad27f92a4d2a922aaa2ccd2f7b30e830393409339232;
// music[7557] = 256'he0311f329337cb36273dd74bb44d4651075720516f4ebb50e84f5050cc4ff151;
// music[7558] = 256'h4956d9527b4f904f234fee4bb045854de154cc4dc94f964d5e494f516b452a37;
// music[7559] = 256'h143eb63e053c993d2a3e2241f4406c419742c73c59398e3923399f366030bb2f;
// music[7560] = 256'h572faf2afd2b072bea2672257c1f8a1a501b161a341427119e12720f1e0bb008;
// music[7561] = 256'h5505f4045e0397fe8ffb9bf99ef5f5f017f2a1f1f6eb32edf0ee0ce9b6e437e3;
// music[7562] = 256'h04e3cbe660e610e06cdfc2def6d90cd91fda9fdcffdb42d996dad2d6e2d393d5;
// music[7563] = 256'h67d315d2d0d0dcd39ad69fd0dcd077d135ceb8cd86cce1dbc3ede6e9b2e8aaeb;
// music[7564] = 256'hd1e7e9e706e94fe5c8ddacd944dba6d90bd945da18d852da48de24dfe6e21ee3;
// music[7565] = 256'h21dfade07ce1c0e0d9dfd2d487ca27cac6cb21ce4ecda6cb2ecb40cab8cf27d2;
// music[7566] = 256'h70d070d31cd349d322d3f1ce1dd2d6d589d278d013d0ffd000d424d3bfd205d7;
// music[7567] = 256'h5fd5c3d45bd92cd924db65dd65dacfd8a8d80fd9cfd6d1d572d8e1d70ed9b5de;
// music[7568] = 256'h67dfb0d7b6d334d760d7f5d9eadfbddfb6dfe3e8adf1eaec67e4f2e03de1e8e4;
// music[7569] = 256'hb5e27ed89bcd8bce7ad940e04fe9b8f1aff2e6f360f54cf5a3f293f2aaf292ed;
// music[7570] = 256'h2deb69eee7fb1a054a00c1002e04a2054d0761082b0c770d670f56117512f716;
// music[7571] = 256'h1d18d217f9186c1cc12111237b251c28f728e52cb232142f0522811f9f21481e;
// music[7572] = 256'h2920d7213d22d1245a26d2260228102e5731752f32302831f6312030df2d0332;
// music[7573] = 256'h923326324a3619366f32b9360c36f83161379d38cc35d137dc372937a639d737;
// music[7574] = 256'hc02e0e2cac3108356635f334ea350632982aad2a842f5c3583332b2e232f1c2f;
// music[7575] = 256'h932f9f2cb428402aa2260426022a2c2e0231fb2bc82bca2c6728eb2716278527;
// music[7576] = 256'h9e258d21d321a21f0d1b2e17cd1703143c0e461d2328561f6c1dd51ea11a8f16;
// music[7577] = 256'h8712c00e830f7b10c30b8f080a069e02e00085fb32fb470021fe79f979f7b6f3;
// music[7578] = 256'h34f1b4f283ecd8df4edaabd8abd7c6d352cfc0d133d2f6d005d1e7cdaacdb2cd;
// music[7579] = 256'h63cb9fccb3cd88cdc9ceabccf5c90acaa5c66ac5c2c86ec7e8c539c72cc8f4ca;
// music[7580] = 256'h7fcdb8cb91cadbccfec97dc7c4cc4ad2a3d6a3d631d760dbf8d72fd6fcd839d8;
// music[7581] = 256'h3fd7d3d6f4d702d72ed671d963d992d866d637d49fd69ed6ccd641da87dd6bdf;
// music[7582] = 256'haedeb0dd65dd55e17ee592e477e65ae72ee5f1e470e257e382e75de75ce7c1eb;
// music[7583] = 256'hfff95a075b03d7fe9b0231042d05e1038e0248062e08e9073907fd05e106bc07;
// music[7584] = 256'hb3073207d3095b10370e0a09530bfa0ae80dbe0d44fb9df494fdddfd0dfd11fc;
// music[7585] = 256'ha5f8e0f418f162f3c9ed71e0d2e1ceec7af2b5f83e01df022b04500222f9a0f7;
// music[7586] = 256'h32f542f1bdf2f2ef28efa0efa6f010f2ffed18ed81eed9f39df6e0f17df60cf7;
// music[7587] = 256'hd6f27af603f8bafb13ff0effd4019503e304d804da088c0ddc0a6a0d88123011;
// music[7588] = 256'h1313db1653160219bc1ec41feb210a25b5241426dc26fa250829bc2b082a7e28;
// music[7589] = 256'h8a29ef2c942e122cac2c822c05317342c149de48a44d784b99471f4a364f8150;
// music[7590] = 256'h794b5f4a174b3249574a544c574c4b4b054b694be7495648e349ab4aad4d7753;
// music[7591] = 256'h3848aa33e92bb82bfb2bcd270328962d9229f127262a562b792ef72ba62b8d2c;
// music[7592] = 256'hb229b22a96297627f023961d301e6a1eba170e147612f10f0d10d40b8a058307;
// music[7593] = 256'h74063900c6fdb6fcc3fbe4f9fcf47eef98eda4eb44e782e4e1df09df82e13ddf;
// music[7594] = 256'h51dda9d93ad8cbd738d187d1c5d546d450d1aad12cd2bdcc0aca94c96aca4ccd;
// music[7595] = 256'h9acb33cd9ccb21c9becd5ccab5c9abc940c400c664c58fc469c43fc8fbd964e0;
// music[7596] = 256'h08dc17e060e273dde8da8bddd6dcc4da1edb2edb97dd44e095e101e092df13e0;
// music[7597] = 256'ha6dc62df35e301e594e5e4dfc1e2d9dea6cce2c994cc46ca3bcc23cf53ce84cc;
// music[7598] = 256'h04ceafcbbdc940cc32cae2cabdcd43d1fad4add1e3d1e6d4dfd354d236d17ad6;
// music[7599] = 256'hf7d83dd5bcd610d7b2d600d88fd521d736da72da24de47dd66d941dce5dbc1d9;
// music[7600] = 256'ha5ddb9dfcbdcbdd969dc7ce141e281ded5d77dd7e2db00dde4e0ede38ce222e6;
// music[7601] = 256'h76ec5bed43ed41edd5e880e7f2e9f6e529daa3d2d5da17e539ea16ee8df01cf7;
// music[7602] = 256'hd5f780fb6f087806aa0b131dcf1dd31b921dd01aba172a172318fe18801de11e;
// music[7603] = 256'h4c1cd31d4d2194254f260e26e2284f2b6a2de82ce5313539f0395c3ddb353026;
// music[7604] = 256'hea27f52bd92ba9319331e1303035e631ed300a37fa37eb36b3377e3c3940403d;
// music[7605] = 256'h463eb3414b43ea448243c544a6459142b342c2445d45f2430244194737465842;
// music[7606] = 256'hf8437e4a164c6647e142c643c545973fcc3cb4424f42b13e6b3dda3ca73da439;
// music[7607] = 256'h2836cd3d7142ae3e1e40aa3d2a37db35052d6427f428b9246f26eb289e2a632f;
// music[7608] = 256'h9f2c2d2d852da328bf28862650266b267a22a320101a331e062f7f2ee5254025;
// music[7609] = 256'hd42416249521011bff153f149f12280f9f0def0d89089f053c06bbff2afe55fd;
// music[7610] = 256'h03f689f422f15af34df878e7f6d808d81dd48dd22dd26fd299d2eccd38cb8bca;
// music[7611] = 256'hcec873c7b8c6fbc55cc44dc79ecce3cbf3c96bc9ebc6bdc73dc99dc65cc660c6;
// music[7612] = 256'h52c564c6d1c5adc671c89ac739c7afc612c627c40ec26cc3b4c3f8c36cc7ebc7;
// music[7613] = 256'h51c5a4c69cc610c2a7c1d1c1c2c019c283c3a6c62fc892c86cc955c8cec983c8;
// music[7614] = 256'habc775cabec775c935cf74d032d148ce46cc4bcec4ce85cd28ce42d170d018d2;
// music[7615] = 256'hf8d4cad0a9d95ce92fea99e906eceaeceaec20ec5cf06ef16cecdcec01f1daf3;
// music[7616] = 256'ha4f1f6edeeeff5f19cf355f562f502f7a6f862fb62fb9ef5e9ed3ee203de20e4;
// music[7617] = 256'hd9e64ee7b4e895ef74f4fded64eb46ea61e60de9f1e69bda1fd3f8da28e412e6;
// music[7618] = 256'h20efc8f7bdf742faf1fc92f90bf491f3b0f311f2b3f1fcedb5ee17f243ee33ed;
// music[7619] = 256'h27ef11f0f1f13cf3f6f3bdf7a4fc2af8c6f659ff86fe54fb43fe0701b004d507;
// music[7620] = 256'h620c560f02100d140d170718a918b7196a1c651dee1e392335246c22b326bb29;
// music[7621] = 256'hed26552a922c962b40313030c72cc131bc3030358547374c9a47be4a624bcb4a;
// music[7622] = 256'he54b554bac4c644c954c404eb94ca84bc648cd457b4518444849044e3e495b48;
// music[7623] = 256'h84499c49d049c53f5e3b0043313f953633368b368a339b329c39223ed93dff3f;
// music[7624] = 256'h8e3fd93e213f763f5e432145af433041d93f6c41b63fbe3a5135e52f912e2930;
// music[7625] = 256'hfe2d2f290226a423542311209f1ae41ac416a71223146d0f170a22054d02d002;
// music[7626] = 256'he1fa2cf8f9f993f338f34df3b2ee77f08eee2de965e956e89de6bae567e359e3;
// music[7627] = 256'h01e1dade04e1d7ddb9d9c2d914d870d785d71fd6f3d691d841d7bdd7abd828d8;
// music[7628] = 256'hb0e311f218f1a9ef6ef2a7ee8aeb4dec91eab3ebb6ee89eddcede3ed99ed94ec;
// music[7629] = 256'hcce9a6ef77ecb3dd34ddafe066e0c7dfece0b6e0cccfbbc666cfb8cc58c98dce;
// music[7630] = 256'hb0cf58cf6cd007cf1ccc6ccbf9cb64cc36cb61ca6ace98d110d4d4d61ed3b0ce;
// music[7631] = 256'h3cd002d397d2b1cf66cf78d223d4d5d3a3d273d276d5e5d3cdd08dd57ed7f8d4;
// music[7632] = 256'hebd600dab1d924d72ad875d883d446d523d93dd8d1d536dae5df77de6fdb9ed8;
// music[7633] = 256'h3bd921dc2adddee25ae43fe219eb3ef0b2eabbe673e4efe318e631e4d9d8d6cb;
// music[7634] = 256'hd5cecfda3adf87e764f055ee9ef23c00460bcc0e4a0cb40a23073207090bb005;
// music[7635] = 256'h8802d90362010f042907250617088109410ab00dfc0eca0fea12de15b419d61c;
// music[7636] = 256'h7319c10ecc08c60c830d770ee813fb1392132e18dd1b1d1bf41b5c1e491e0824;
// music[7637] = 256'hdf2599238a2cec2f7d2b272d732f713065302a3220344333c234ca3414347236;
// music[7638] = 256'h5d3533347f36bb3463301d303f3109338c36eb38bd3906374630302d22306a33;
// music[7639] = 256'hdd350d370d35e1326530902c092a562d2335af3643347e339e30922d0c29d326;
// music[7640] = 256'h282b532cde286a298b2d202f9d30a02f0e2b7e2bde29202758262c25fe30543b;
// music[7641] = 256'h9d388837a932f52c4e2cb4278d232a24a121f61c9b1e0f1e6d189716a312c40e;
// music[7642] = 256'h20117d0eac0745079d060904fa0442fa7fe740e20be3acdfa3ddeedc0dd91fd8;
// music[7643] = 256'hb6d95dd590d46ad24dcc8ccea7cdfdca43cf9cd112d192ce2acddfccc6cd8fcd;
// music[7644] = 256'hc3c899c98ecba8c748c5efc3aec44fc49fc1b1c38bc674c5cac491c34ec26dc8;
// music[7645] = 256'hbfca5ac59ac7fac7abc22fc39fc97dd419da17d93cd93ed9b7d90ada97da29dd;
// music[7646] = 256'h77dfedde04ddb6dde7dcb7db6bdd5cddfdddcbe04de41be6f5e26ae023e17de4;
// music[7647] = 256'h11e6cae473e7c5e43fe53ef793ffc7fc47ff39fe95ffb6016900460181fd93fe;
// music[7648] = 256'hdc02b8fffa007d01aaff9b036005b304fc043b0462048a0504042805030388f5;
// music[7649] = 256'h01f49af745ecdbe88beee8f1f0f5dcf7d1f7a8f81b00c80472fd21fb41fceaf8;
// music[7650] = 256'h40fc1bf922e6dce451f1f0f3f0fb3cff47fe060977090a08fd0786fb9ff406f1;
// music[7651] = 256'h96ed3cf0a3ef35effbf1f7f282efb6ebafec85efa0f0beeff5f0d7f2b7f579fc;
// music[7652] = 256'h71fdccfcf8024b06e90446057309650e4b0e8c0e5f125f11ad13021ba61aee1a;
// music[7653] = 256'h061d9c1faf23a61f7d20ea240b2461273328b527d825e229703fd24872454246;
// music[7654] = 256'hd7424143e2453a46904b7e4db54bc44a5a472247914c254f984db948c646954b;
// music[7655] = 256'h26484242cf46b44a304da047c9354c2e0b31e22c3f2be43244357531882e942b;
// music[7656] = 256'h6a2b58282a2408275526d1246d29042ade28d32a472bdb2a442a69270e27f029;
// music[7657] = 256'he5268121ea21691f2b19e2178715b21123121e10fe0c1c0b1405bf009500baff;
// music[7658] = 256'h41fe78fa82f4cdf047f03deef7e90ee879e60ee582e755e606e1e4e02cdfb8da;
// music[7659] = 256'h7adcacddf9dbb3d92bd78ed92ed76ed018d293d1b2cc35cd92cf38cf5eca20c9;
// music[7660] = 256'haacc27c9c6ca53d80ddecadc9fdfd1e0b1dd8ddc8bdd87db94d927dc1ee0bcdf;
// music[7661] = 256'h78dc50dda3dcdbd855d84cd903dd5fdd9bdbdddd72db95db2fd64cc691c4bdc6;
// music[7662] = 256'hd7c5f2c77ac5d6c7aec92fc8adc923c69ec81bd07ecd94cadecb24ce00d138cf;
// music[7663] = 256'h6acdfbd152d3a2d2d4d485d4d0d543d551d256d473d557d768d752d660d9c2d7;
// music[7664] = 256'h6fd76bd84ed79ad99ad8c1d863d92ad779d802d80edaf6db0dd93bddd6de87d8;
// music[7665] = 256'h3cdbefe0b7dfabe203e3b2d9a2da50e06fdf37e4aee889e58ce7cfeef1ee42ea;
// music[7666] = 256'hcde7b9e40ce14de1dbe299d661cbf4d411db52e5ebfd2607420a9f11ea121210;
// music[7667] = 256'h6411431e2d23b01afc19711c711a4a198c1a881a1b1ab31cf01fbc20001fae22;
// music[7668] = 256'hf02535248e28ee222c1361121919f01b251d381fe221d5244c260226932c6632;
// music[7669] = 256'hd4302b31ab31e8345238f935de359638843b3a3e943fd03eb63cdd406345fe43;
// music[7670] = 256'h6146f7477a42e9413e452447584ab1476243ef43b543a446d3479e476a4ac345;
// music[7671] = 256'h26448848f644f740f740d1418643a74486446544b2444241dd3c383e2f440746;
// music[7672] = 256'h4042fa42f341ae3cce3c8d3b4a37fc30e1298c29752c572cd527f728cf2baf23;
// music[7673] = 256'h632a7b3dee3c95360938933885359e31f12fd02c362a5129cb25a8230122df1d;
// music[7674] = 256'had1911159c11840f220c860ac00a7e06f2047b059cf526e62ce764e41be168e2;
// music[7675] = 256'h27de98db97d98fd64ad8b2d870d758d760d621d471d23dd367d185cdb6cd9bcc;
// music[7676] = 256'hf0c9e2cb51cd3acc65cb74c6d6c3bac71cc685c206c487c420c6e1c8f3c6d1c4;
// music[7677] = 256'hbdc5a2c3fcc1fbc50cc61fc0c2bcdbbf05c45ec064be59c2f9c1a3c283c440c3;
// music[7678] = 256'h8fc4c9c4ddc3d8c4b4c3dbc289c189c012c5b8c696c581c759c648c531c590c4;
// music[7679] = 256'hc6c826cc25cc37ca8ec944cca8ca6fd1d5e2dfe85be8cde916ebd1eb84e921e9;
// music[7680] = 256'h9bea2eea99eabcecedecf7eb87eff5f056edd7edb6efe4ef19f1f1f075eeebf1;
// music[7681] = 256'h34f471e5ecd8f5d96adad1dce5dfe1e059df9fdb6cde2ee03ae050e54ae6c7e6;
// music[7682] = 256'hfdec0bf3b2f259ed33ea80e819eaeaea50dec5d195d738e1b0e308eb1ef250f2;
// music[7683] = 256'h3cf796f981f4d4f3c9f3aaf0eff075f0f3eccbed1ceffeecfcec24ed2fee4ff0;
// music[7684] = 256'hbaf01ef36df51ff65df7b1f888fbb1fdb3fe59017903a3046408fb0a370dd612;
// music[7685] = 256'h39139413fd175017851aad1ecc1e0e221d2279223a2442251e289b26dc2e9040;
// music[7686] = 256'h6745c544df45dd449e4449464748294a0c4b6d49604a484da94c1d4c1d4cd94b;
// music[7687] = 256'h894ad44b784f2a4d424b944ac849f4474138ee2de031942f292f3e30c62bc02b;
// music[7688] = 256'h502dd73063364134522f762fc02e702b782dff2ede2b4832f83dbe3f993e1640;
// music[7689] = 256'h7a3f133f6e3f6d3faf40363e263a843b273b1c363e336f312a2f6a2d6c29a525;
// music[7690] = 256'h7e23731e4c1a99185f15b5128b10bc0dc709d605fa05e304f9005400a6ff48fd;
// music[7691] = 256'hfbfb6ff913f638f4a4f2f5f03aeedeeb91ecf8ea3ce92be97ae48ee3e7e3c6df;
// music[7692] = 256'heedf8adc7dda74deb5dc0ee623f5b6f30df121f2b4ef03ef9df04ff041ef89f1;
// music[7693] = 256'h4cf150ee5feeb3ed6aed0fef9eeea0ec86ec83edeeed20efa0ed7aef1cf085df;
// music[7694] = 256'h4cd556d516ca51c4f0c531c4f3c4f2c576c733c7f0c42cc51ac5d5c6e4c96dcb;
// music[7695] = 256'hc7cb61cb3bcdffcd47ce2fd0cace6dcef0d00bd082cec0cfb8d0b2d03dd018cf;
// music[7696] = 256'ha8cfa8d02fd036d182d383d694d750d372d085d14bd2a0d474d690d4f8d31ad6;
// music[7697] = 256'h4fd8c0da56dc0fdbfed946dc27ddbddc90deebdf09e2c4de08d672d807de2bde;
// music[7698] = 256'hf1e1e8e3e7e248e779eea0eda6e74be79ee37ae258e75bdedfdaeae914f2f4f4;
// music[7699] = 256'hd6fb6301bf05ad09d40ab40a4b0b970a020981062105c805ae0211004400e7ff;
// music[7700] = 256'h51005901cc03cb038706b40810fa84f1bef761f836fc8d00e0ffa1032d054e05;
// music[7701] = 256'h2009670c790f26127215e2198f1b1d1ba41c471feb2120244024a0256328d229;
// music[7702] = 256'h812a9d29822b672e102d4a2e262f742cfa2f1b3469318e3166347d32e3304f32;
// music[7703] = 256'hfb320e33f632a4339a357e366e35ce34bf349b332b334f328a326737c338ea35;
// music[7704] = 256'he8347332992f692e9b2e7f343d3948348f30852ff829482a862bd627ae29242a;
// music[7705] = 256'hd82a3f2d182cc837dd45714537437041813f5a3eec3bdb39f537bd36ea33da30;
// music[7706] = 256'hed2d492966279724d620941f6e1c4f184017f4159c104c10050d68f9e5ed8cec;
// music[7707] = 256'hefe74de9e0e718e325e368e059de73dd95db5edbc1d9c1d89fd869d748d76cd5;
// music[7708] = 256'h0bd3e5d314d40dd357d138ce14cef2cde7cba9cc3ccbd6c751c95ecb10caeec9;
// music[7709] = 256'h4fcbefca39ca10c83cc692c640c431c4bdc51dc4f6c54bc721c68dc788c7bac6;
// music[7710] = 256'h8bc7e4c72ac87bc8dec654ca7bd676dc92da2cdb35dc37dc95db67db5bdb77db;
// music[7711] = 256'h6fde0ee09be041e1b6dfd5de3fdefcdf31e1f1e1ebed19fa43facbf86af823f7;
// music[7712] = 256'h61f8f7fa8efb6dfcbcfce7fa09fd6cfe45fc9bfd5dfdc6fb1afe6e00e9000200;
// music[7713] = 256'h24006e01300379fef2ee52e8b5eb27ecf0ee69eeaeec77ef63f025f4cbf17de9;
// music[7714] = 256'h94ed66f484f5a9f8cefc37fdccfdee0257047e010aff31fbdaf972fbdff70deb;
// music[7715] = 256'he7e381eb1df260f78cff95046d08890a690cd00bee06d304aefe16f437ef27ed;
// music[7716] = 256'h26ebb7e90ceafdea4eeafdebdcee0ef041f26cf589f81efa2ffa95fb8efec001;
// music[7717] = 256'h4103c603aa05a008640c140e0c0f49124d13161477168e195e1d171da41e7820;
// music[7718] = 256'h512175302c3e583cb93bbb3ddf3f574228438645c846d4468347c84657476f48;
// music[7719] = 256'h57470847d0476f4713471a468145ea455847fa4ba8451733072dc72e622c6a2e;
// music[7720] = 256'h0c322c327030bd2dfa2baf2a24292a2afa3050369633f831f332002f982aef29;
// music[7721] = 256'h072a492bd92ca82b2a2bad2de82df32af529ec2ae82af42880254a245724b121;
// music[7722] = 256'h1d1f351d2219df1487132211bf0b480aa80811036001fc0062feb2fb7bf98ff7;
// music[7723] = 256'h9df286ef4defa2ec2deb6fe963e680e483e1fcdff1dff8dd7fdb19da6fd7b7d3;
// music[7724] = 256'h04d25fd1efd25fd247ce87ce09cc75cd48dd34e553e234e2f1e031df27dfddde;
// music[7725] = 256'h96df15e02ade94dc2dddb8dcd5db40dc7adc80db6ddc70de86dc5edcf0db1bd9;
// music[7726] = 256'hfddc34d785c62fc49bc815c83ac7acc5ecc482c64bc771c637c85dca8ac945ca;
// music[7727] = 256'hdacb3ccd60cf6ad0e6d0fcd047d077cf15d078d147d123d1c7d040cfffce49d0;
// music[7728] = 256'h05d101d1bcd13ad3a2d33dd288d21ad4c1d3a4d46fd414d36fd3fad0e0d03cd4;
// music[7729] = 256'h57d4ded4aed533d620d820d9dbd9b5dac1da6ddae7da58dcdbdc1bddcddd45de;
// music[7730] = 256'hd3df8ee080dbf8d865de2ce078e116e6c1e4bae52fed57f10aefc5e8e6e91df5;
// music[7731] = 256'h95fdfbfbe4ef79e6b7ec8ef580f9720110082c0aa90d500ecf0cc10c02097307;
// music[7732] = 256'h7b0f7816ac15ad13f0138814731560172b1263079606f509260aa00c510d5e0e;
// music[7733] = 256'h0111b5124b17ed19f31a3f1dca1e7c2103239726cb2c202f9c300f314831d533;
// music[7734] = 256'hd434fb3599370a37a137e739293b1a3c153eab3f3940c73fa53f364116429a42;
// music[7735] = 256'h71435b43be447e442f41dc41334484445645bc441b4491464d4817470846a545;
// music[7736] = 256'he8435b423342bb44ee4734467644904361404d3ede3c46417e4792440a410c40;
// music[7737] = 256'h573eff3b763b633c3039543f764aed446c3fd04172411841623f903c813b6a3a;
// music[7738] = 256'h49383436ae34d031612fea2cef296827fe23ab21ca1e331c671a70176116190d;
// music[7739] = 256'heafd25fa74f801f4f3f277efc2eb2bebc8e921e807e621e40de3bbe035dfa5dd;
// music[7740] = 256'hc8db1cdf6ee138dd03daa4d84fd64dd466d27ad0dbcd80cb2dcbdcc903c87cc8;
// music[7741] = 256'hf8c665c4a0c439c4d0c3ebc353c3f7c34dc3fcc27ec3e1bfebbc89bd25be95be;
// music[7742] = 256'h2fbf07c03ac046c01ac173c190c108c27ac275c2eec2f2c374c465c565c5bdc4;
// music[7743] = 256'h5fc5d2c593c6adc683c686c7a9c73ec85ac8c0c861ca22c902cf43dd9ce240e1;
// music[7744] = 256'h4de2f2e2f4e233e4f4e4dbe4b1e5eee5d9e58ee689e6d9e634e719e83fe922e9;
// music[7745] = 256'hd9e917ea59ea59ea16ea3bec0ae5c2d7b6d5a9d7ead7a3d9dfda3fdd00dfc7de;
// music[7746] = 256'hf4de73df8fe04de357e5a6e043db1cdf82e4efe7c9ec2eedd2ebf6f00cf642f3;
// music[7747] = 256'h77edd0e9d8e6e4e639e9fce0c7d274d4e3deb1e22ae9f1f070f3c0f7a7f959f8;
// music[7748] = 256'h00faf5f8d2f5a9f309f1d2ef27ef06ef33ef83efc7f08df1b6f290f326f6ebf8;
// music[7749] = 256'heef4bdf297f526f7b7f9b8fb2afd4dff9900ca024c0498067909bd0ac20da80f;
// music[7750] = 256'he011bb14da139a1c962c7e303930513311348735b437593876395f3ac33a963b;
// music[7751] = 256'h523cc33c6d3db53d8c3d083edc3e583f963f4d40ef3f1f40a1401637fe2c252f;
// music[7752] = 256'h132f752ce82db82c052b7e29982a242f472e762c082de82a91283f260628ff30;
// music[7753] = 256'h0533062e582f492e122ac22acb275926e8266424cb3258466d4660445146dc44;
// music[7754] = 256'h2446ea47dc466e45d2431242e43f463e943b6836bc321b30822c392918278d25;
// music[7755] = 256'ha722f01fe91d1b1b9e188e1518139e104c0dc10b4909aa060205a002660171ff;
// music[7756] = 256'hfbfc49fae3f764f743f595f346f12ceffceec9ebd8f2e200670133fed0fd2dfc;
// music[7757] = 256'h12fb47fafdf9f9f8ebf7c5f69af5c6f5dcf4b4f44ff447f34df36ef2f7f195f1;
// music[7758] = 256'hd8f128f1e9f0fef175e87ede37de43ddd4de15e0abdf70e0cadea9df57de5fdf;
// music[7759] = 256'h1de087cce2be43c30bc2cfc2c9c525c32bc3c3c364c4c8c6c0c64dc53ac426c4;
// music[7760] = 256'h74c5a3c5ffc406c609c707c7bac7b8c802caf9ca07cbc6cb01cc80cc79ce3bce;
// music[7761] = 256'hecccf5cc46cd2ececdcd67cd00cf17cf85cfa6d049d167d4a4d50bd547d65fd6;
// music[7762] = 256'h59d640d67ad5c8d51dd604d736d96edbc3d7d1d015d221d705d9d1da4addb5dc;
// music[7763] = 256'hc9dea0f07fff3afb38f7e9f42ff196f394eed5df5edd07e78aeb8bf0bdf848fb;
// music[7764] = 256'h3efe370089ffbd0056ffe7fd75fdebfb4bfa54f947f8c7ed43e366e59ce88fe9;
// music[7765] = 256'hcaeaf7eb05ee23ef20f158f3d6f580f81bfab2fcb3fe7f01fc055e09230c910d;
// music[7766] = 256'h3210d1133f167519431aa519221b7a1bf51b121e8b1fc5204222fd236d25bd26;
// music[7767] = 256'h8e28e32740264827df28b62aca2a5829e62a1f2c1a2d6c2e172d2b2d312ef32d;
// music[7768] = 256'h902d272e7e312b3205307d2fca2d532c232bc3298d2cee2e922db42d1c2df029;
// music[7769] = 256'h1e28df286b2f6433b52de92cd22b3c27b931533da73c703ce63cb83c823d883d;
// music[7770] = 256'h043de63bf93ade392e38aa36023525333631e92ece2bc829802792249b229e1e;
// music[7771] = 256'h1c1ddf19490b9f01ce01befe43fbbdf8c4f527f451f16fee23ece0e927e875e5;
// music[7772] = 256'h56e39ce1cedf68df96ded8dcb0da65d94fd84bd68cd6b4d52ed1f9cdd0cc88cc;
// music[7773] = 256'h74cb16ca9cc950c89cc738c734c6cac52ac5b7c456c429c4d6c3f0c1ecc0eac0;
// music[7774] = 256'h73c06cc079c0e4c08bc06bbf17c068c0f6bf26c2d8c42dc5b5c591c68dc51cc6;
// music[7775] = 256'h2dc65ac5fdc7c8c5a8ca8ae0bbe930e708e99ee8b5ea74ecd2eb31ecccebedf6;
// music[7776] = 256'h450327027e01320312034203490396034b04c4040d0456048d04f2034405bd05;
// music[7777] = 256'h03067706b30688070e072d07870765093d099eff50f9bdfaa6fa5bfa9dfabefa;
// music[7778] = 256'h05fb76fb1dfc1ffc10fd80fd93fdb0fe50ffa4013406f0051aff0dfdeb012b04;
// music[7779] = 256'ha906d8094207f2068f0ee8111d0d9b091b07de03f105300569f762f027f952fc;
// music[7780] = 256'hd4fe4108df0be20d4c0feb0e7f10f90f200e150d920d3d01d1e999e40ae7a5e4;
// music[7781] = 256'hc4e4f4e211e40de662e62be976ead0ec05ef8bf160f4abf577f80dfa09fdadff;
// music[7782] = 256'h5500b903f604b3083c0b1b0ca01afe26d526bd285f2bec2c802fa1302f323334;
// music[7783] = 256'hd634bc3575360c37f3377e39bc3cbb3dbd3cf93c893eb742b3438642b4446346;
// music[7784] = 256'hb448e149de4767463246ff48c94aeb488a47ef46c0455a43c34224452b472d47;
// music[7785] = 256'h30485a4ade45f0414f43353c7b31212b79261224942171204d20b71ef51e2b1f;
// music[7786] = 256'h2d1ff11f591f4d1f0a20fb1fb81fe51e011e731c5519f216d2146212cf107b0e;
// music[7787] = 256'h8f0d060cfd061103fafdcef9b7fa68f9e2f5b0f29aefc9ec31e8f3e785ec97ec;
// music[7788] = 256'h29ea8de664dfbadb05da52d59cd7fadfa9e27fdd8ad42dd099ccb0c537c4e8c5;
// music[7789] = 256'h2ccacfcee7cdc1cee6ca8fc287c118c066c010c208bf60c2b1c572c377c359bf;
// music[7790] = 256'h4fbbb6bc9dbb5abf6ac877c56abc5dbd3dc11fc16ec070be6bbcdcbb3abf97c6;
// music[7791] = 256'h23c80ac889cbacc8b0c3e5be0fbb93c2a7c921cd78d387d1b6cecbcbc2c30fc6;
// music[7792] = 256'h11cd37d547ddfcd6e8cefec910c672c96bc796c62eceefcc20c83cccb5d624da;
// music[7793] = 256'h71d044cbe8ce73cffcce2bd570dcd7d9f8d0d7c72fc3ebc69bcc5ed55edecae1;
// music[7794] = 256'h71e213db6fd5c8d8c5d9a3d9f4d84add45e0bed45ed4d6df98e3c1e224dad7e1;
// music[7795] = 256'h5cfdafff78f8e006e413ca129f0ba806710857098e0db21b15214218a11a8a2a;
// music[7796] = 256'h852a8e1cb71e3f2e82375e379932242c3c2c963935420b3e66374130a037d848;
// music[7797] = 256'h5a530458264c2f42274c3451144f274e2c4ef055505d2554dc4bdd5b52663758;
// music[7798] = 256'h0f526d66d178f666a44df44baa499242dd4398468346264c1d500f4c4249e741;
// music[7799] = 256'h8047f55efa5f1e506c47144de151ce43f03ce444174e705570527b42272b3e26;
// music[7800] = 256'hf931693b85406b31021fab27c93b1b3bc42759195e08a309b1225628dc22d11c;
// music[7801] = 256'h101c7a1b0e0363fa380b0f13610fb7fee1f55502aa074df9c7f11ffd1204cb00;
// music[7802] = 256'hd6fa35f722fb6af54ce473e163edc9f237ebe8e0a5e427ef10effcee88ef72ed;
// music[7803] = 256'hfced0beddfeefde68ae062ee50f505eaa3c8c4af9ebd96c1febbe1c6abdabef5;
// music[7804] = 256'hfef55cd373b30aab02c250e115ee38fa4110240c51e8c9c993c141cea5e0e6eb;
// music[7805] = 256'hdceaa5e256eec900f5f98bec19f41d09ca187f25b129b016d90304066609a20c;
// music[7806] = 256'hab17010cf1f6cefae0fc0c00550f8c15951afc1831095202b408160e7b076df9;
// music[7807] = 256'he2f0e2f024f96207fc13c9251739c4310b187d08cb0da41dd71bc018e0221029;
// music[7808] = 256'h4b312338e53f074c1e4efa498d372923312c623f523b56288f2954393537f42d;
// music[7809] = 256'h57326e3a32318219150319f635f81401fc06700be20e690c870059f8b0f4f4e5;
// music[7810] = 256'h9ad853de64e8bfe826e61ae23ee285eabee473dbe9eb2df8caef16eb69e56ee7;
// music[7811] = 256'hb0ef0cdd70c6b9bb5cb64bc74ad43cd6afe4bcebdee192d404cdbcca46ce25d8;
// music[7812] = 256'h60dca4dca4db19e2ede9d9da26da7cf019f4c6ec9fe37ddf35e41de315e9abf3;
// music[7813] = 256'hdcef99e8d8e862e8aee43be955f0f3eef1f4c8034203a1f543f6bcff2ffb58f5;
// music[7814] = 256'h55f3edf016053f19d10b49fbbbf967006306f6027f023502c4039c0e2016271f;
// music[7815] = 256'h5c1d3c0787fadaf8c3ff2d112817e6159c1b8c1f0d25b82f5c3069271a237e21;
// music[7816] = 256'h351ffd1fa41dec14e50ed2080508e913f11628173e249826a41d1b180917a61f;
// music[7817] = 256'h2c2814283c2a3b2cfd25541fb51d8919930ff513b12a822d571edb19401cf827;
// music[7818] = 256'hfa2d9222f0185a0e39117d22751d6013e516e10cacf523f1c9feddfbadefb7f3;
// music[7819] = 256'hcaf78afdd70945017bf5e6fb93f8caf7cb0b7b13a00a870723097f06cdfbe2f6;
// music[7820] = 256'hac03ff07d3f511e8c3e449ebf4fa10f7cbecbeeda0e785f145048a0094004201;
// music[7821] = 256'hc5f5c7f35ef505f2fef213f7c2f687f454eef2de3ddc6fe80df1f1f787f509eb;
// music[7822] = 256'hbfe39ae336edfeeafdddf2db46e1c2ec15f75bf5aae7d8d718d982e6dbedc1ea;
// music[7823] = 256'h0bed26f90cf481e7eae2a4dcafe782fdf50094f67ee934e32ce4bce824ed96e8;
// music[7824] = 256'h57e6d0ebf5e569d277c6f8cafed2d7d9b6ddb1e0e7edc8fae6fde5f10ddbfdd5;
// music[7825] = 256'h70d1b8c05ec5d5d2abd9d6e0a0e19ce14ddf20ddcae3b6e6cee6dbe783e3e5de;
// music[7826] = 256'h87dbced6dcd9bfeddbfe72fd9c018b0b56ff18edc9efe8f8dcf9f5fc8703e606;
// music[7827] = 256'h810bb1123619311c3e16dc0df410a71b8b22e128c02cb928132afe29d91f8122;
// music[7828] = 256'he52a562e1338ce3c88384b311e30d436c833c034ba3b0a3b12418041573acc39;
// music[7829] = 256'h9d36163bb3413c3d3f3cd63b06397c3cf13ed338b8325f370442d9440c39962c;
// music[7830] = 256'hb12bf72d9d314a33bc3026351636b72ba3265628342b912f1d315f2f9b304432;
// music[7831] = 256'hbc269619f121f22dc4294a22ba1d5e19651897162715f11b591b37111c10d50f;
// music[7832] = 256'h140d3911c713200d39058408e60e2e0b72003103dc11630b3003f604fbfe6f08;
// music[7833] = 256'h9d07aef870fe00ff6d037b0a09029dfc80f195f862121713780c7e08b1021f01;
// music[7834] = 256'h1afe04ff31048b06160232f8b7f1caf1b2f815fd4bf744f0c0ec13e7c6e2a1e6;
// music[7835] = 256'h62edf0eed5e83bdc6fd23adb6de8b9e3bce4ede819e228e3e4db83d3b3dd77de;
// music[7836] = 256'h14dd9cd802ccc9d9afe2efce34cc70d391d78ce153dd8cd26ec9a8bbd2b317ae;
// music[7837] = 256'h67b406c1efc33fc714bf88b6e2b8a7b4deb60ebb75b93aba13bc21be3abb95bb;
// music[7838] = 256'h39c17fc235bf8bbd57c10dbcdfbeecca81c2cfbe62c2bec090c0beb852bca5c8;
// music[7839] = 256'hb4ca5fcc77cbdbcac2c8c7c357c482c3d6c6fdd184d8e7d892d1aac88acc4ad5;
// music[7840] = 256'h3cd620d7dbd9a2d638d2eed35ed721dadadcc4d73ecd46cb7dd569e293e6d2e5;
// music[7841] = 256'h63e404e853f6c7fbacf88affbc04800119ff6102da0d3316990de304c50499ff;
// music[7842] = 256'h8400320ad5117019bf160413fa1b78236b21ce174a123615e6169119c31d6623;
// music[7843] = 256'h53285b1fbf12571ab027a12a672a8e26b4283e316a30e92b70272f27f429372b;
// music[7844] = 256'h46329933a128371ca322bf3708355730a636762c1f2c69338d302133f630e52f;
// music[7845] = 256'hb4371d33fd29df2cab31a53281362635522c222d9e3586386e39ca35bc2bc22f;
// music[7846] = 256'hbd3cfa3cbe3a7e3cac41273a31298c401c54163dfb40074c06433f4a54458d37;
// music[7847] = 256'h1d3b283aa83b704378432d469f48b740f53cbd423e47a047a8411a3bc63d2149;
// music[7848] = 256'hc54d40408038a63ebb3e903ec2459b4baa4820487c47d23d2b4282482a43333e;
// music[7849] = 256'hc82f412e0d3c6c3ef73aee35d3373236353238381a27c910d415d41deb1f151e;
// music[7850] = 256'h6a186e0fde09ba0a63062905100bcf0f9b0ec5069808090b700836102f0e6500;
// music[7851] = 256'ha5fb8ef82bfcd90608057b010f08ab0b090a490477fda1fe6cfd48f689f9cc05;
// music[7852] = 256'hdd099a01d6fbb3fbdcfacdfffc01b4fc93fa44f58fefe9ee4df50c06de0ab502;
// music[7853] = 256'hb7f81bedd3f44cfde7f4f6f7bafbf4f8a5fa33f3e6eefaf371f1c5f24af94bf7;
// music[7854] = 256'h61f51df64df698f4eeed55ee10f1dae9e6e96cf087ed17e7fbe527e9ece97ae8;
// music[7855] = 256'hbce98ae985e64ee69de6cee227dedadc89e32ae77ddfa4dffee1a4dbbdde6ce5;
// music[7856] = 256'h2de233da59d43ad73ddd97daf8d4b4d717d9c5d304d53bda0edc8fd702ccbcc6;
// music[7857] = 256'h4ac9d4ca96cf27d560d16ecdf6d016d1b6cfbed14bd270d0f9cbc6c9d9c6cec1;
// music[7858] = 256'h9ac4b6c9e8cbc7cc2cd262dbe5d070c1c5c6c8c931c590c5eac4afc3bacb01da;
// music[7859] = 256'h61d8ffcdbacda1c952cd43dfeae5e7eafeeeede5a6e0cbddfcdbc9e3c7e4fcdd;
// music[7860] = 256'h8edcfbdef4e341e2e4ddb5de5dd6a2d46ade22da31dbc3e6cce6c7e148db56d4;
// music[7861] = 256'h9dd2bcd53edac9dcf4deafddd0d915d9f7da4fdaf8d807db5cd5a5d310dd30d8;
// music[7862] = 256'h2ad0f8d3e7d6e3d68ed55ad481d8a0e22cdb19c5cdbb07b58fbcfed2b1d5bdd5;
// music[7863] = 256'h09db34dbc0dec5dac7ce11cfa8d5f9d035d4dce414e14ad683d6a7d113d14ad7;
// music[7864] = 256'hedd9f6d989d82cde8de1fbd8c3d48bd803de61deafda8fdd5ee019e1c2df31dd;
// music[7865] = 256'h38e006e0c2e018e4a3e7ccee71e833e4ede5acdfffe767eee4eb7cf306f219ef;
// music[7866] = 256'h76f343ebe6e0d3eaf3f4e2f3e4fb27fe8ffdab0490fa59f298f393f061f67bfd;
// music[7867] = 256'h230096ff3ffbe1f8a7f7c2f780f8eafefa05db028bfd18fdb404ef0429fb7dfd;
// music[7868] = 256'h4f022b0442051cfca4fa3eff22f463ea78edabefc4f1c6f519f538f1e0f46dfc;
// music[7869] = 256'h66f76af2aff779f935fddd00910033044703abff95fcfaf605f92903940ca307;
// music[7870] = 256'hbdfa31fd8201cdfe04038d05d606790e5c0f5d076b021f06590c450d5e0c250b;
// music[7871] = 256'he90cc70fff098a08b30f8311bc101a0f690f6214d118f11fdb22a018ed136f1f;
// music[7872] = 256'h2f2208162e1c7634f84129410d381932f834ef36fa3de94736430a3c87407e44;
// music[7873] = 256'h4443cd3f5738a137b8421b4827450745eb43723c0c3aac4474484145414a0844;
// music[7874] = 256'h8b3fc549d3464147ce4eef4b924bbc464b44e9471f4159412b497d4a6c494b48;
// music[7875] = 256'hda479b45ee450e469a4530440a2f9f238a311530ec2bda2e08278c2494231222;
// music[7876] = 256'h9c2acf2d2c2f39328d28c21b2a1c2727252d842b072d572f842d5e274a203a20;
// music[7877] = 256'ha7259825d5226c27fe28b427ae29ac1f43141b1b4228a82836241d2dfc2da228;
// music[7878] = 256'h022f232ba0274428cc2007252229bd2957301c303d2e7e2966244926fc229c22;
// music[7879] = 256'he52816281e2461278a2eb22c57253825962599254a2a67281c21441f79226325;
// music[7880] = 256'h8322e623a327aa20461b37208a28f2268a224525b11bf0176720001f5123de20;
// music[7881] = 256'he21647181716df16c817ab135014f010ec0f4811310f390df30b700eae0b9d04;
// music[7882] = 256'hd405940c4b0d25064807f40cd90dd608c0003b02bbffc4f949fda3fa90fcec00;
// music[7883] = 256'h68f70ff7ccfb18f147ec3bf261f0c9f0f3ef2ce504e9a2f163ed7ceba3eadee7;
// music[7884] = 256'hb2e841ea4de6dde1eee538e4c8dd3ae825f788f6a3ef09ecdde9afeca4ee24ec;
// music[7885] = 256'hfcf54a0a0114de0b10fe43fa12fe58019303b604bb021401fd02740207fff4fb;
// music[7886] = 256'h45fa59fb18fa9ef76bf941fb29f82df6bef6b3f2eff1aef536f28eee02f2f5f7;
// music[7887] = 256'he9f7f4eed5e94cee61eff0eaf9eb89efd9f01bf28def62eb60e9eae8dce9b5ec;
// music[7888] = 256'h66ee41ec68eb5ee3e1d2e1ca49c599c218c814ccc5cd83ca44c62cc842c8d0c5;
// music[7889] = 256'h0dc519c640c5a6bdffb9aec26dc20dbc76c3b0c32fbf65c124b8ccb0f5ae0ba9;
// music[7890] = 256'h00a41a9d39a0daa65ca0e49aff9b1e9d1f9f3ea4dfa40aa3f3a3249d609a87a2;
// music[7891] = 256'hdea60fa2df9bfea1f7a2949ad6a2acaa1ca491a01ea6b7a98ca4d49fb29f68a6;
// music[7892] = 256'h54aed6adf5ad91adabac07b09bb25cb25eaf45b1fbb276b0afb2cfaf0aace3b0;
// music[7893] = 256'haab983bf74ba1bbb59bcc6b6f2bfeec225bf1ac5a2befebb92c23ebfa5bff9be;
// music[7894] = 256'hf9be30c8e8c5eac177c7a9c676c6f9cad6c904c6efc6e8cccacdc0ca8ecb78cd;
// music[7895] = 256'h66d23fd280c928c912d08cd3e3d224d38cd451d2aacd31cef1da2bdf2dd7d8dc;
// music[7896] = 256'hdcdf54deafe123dc37dd58e0eedec6e5c1e549e3e8e6a2e50ae2b3e488ec2eeb;
// music[7897] = 256'h0ce62aeaa6ed99e890e77bf257f575ef97f20af78bf812f8c5f530f96509f113;
// music[7898] = 256'h1d0d4311b21bd91ef021e6193c174d1dd420a8269a21a91eaf256d220f1c3f20;
// music[7899] = 256'h0a291525ec201b28ba291529732c4f2eb32899257e2c482a7929aa33db33ec2e;
// music[7900] = 256'h2533de3702340c353f3aa639653b033a7b34f23317388b3d9443e84c3b47a13d;
// music[7901] = 256'hc345213d8c2a242f7433663002334f310c2df72f5531c031b434c0372e3bfd35;
// music[7902] = 256'ha534993fd140d6411547de3f013b3840bd4320451043073fc141e847d845ad3f;
// music[7903] = 256'h0b447a4ca5493a44aa469f4ecd4fcd48a54b284e6c471249414d964dca4ef34e;
// music[7904] = 256'hab4c904b834d704d214f2a52954f584d694d274e2850b956cf55ad4cca503955;
// music[7905] = 256'h1158b85d0d53cb4a7250ca571d589f55135d155cdb55cc543c51845565517349;
// music[7906] = 256'hed53f560c26ab069a163be64775e9b584a5d1463536483633f673b65465b5f58;
// music[7907] = 256'h2b5c135fee5e8b5ec15e12585a514d54eb55cc56575cc45b2e59a956534ce449;
// music[7908] = 256'h1356fc57264bd646a84d114fb149ef498f4df94bc04b32471740f442e040563d;
// music[7909] = 256'h8240963e723f2140273d9c3c16357b2cd52d61358b3b0c3b4638cc33f92e392d;
// music[7910] = 256'he92aca2a3e2f2831ce2d0f270c20f51e4f24cb262522eb244034b636012e1634;
// music[7911] = 256'hcb3ee63b6b34da38e53b3f33063720368f21bb1abd198f121d14f916c5174217;
// music[7912] = 256'h4312c30fd50f040f7d10bf127a11bf106c0fd90ab80cbe0c640332fdf2f94d01;
// music[7913] = 256'hf50ba104f702a306c901d003c9fedaf7f0fd20fafaf0dcf30ffbe3fb2cf85bec;
// music[7914] = 256'h46daa5d637da12da22d676ceded25bd680d47fd408c9b9c35ac68ac37fc3f5c6;
// music[7915] = 256'h0bc96ec138b9a3b918c080c6e6be4abbd1bad3b367b757b94ab8cdb462ab1eae;
// music[7916] = 256'h85af7daf0db34ba9d09e3c9d5b9e0ba0a39fe09f55a061a0cba0e39d4e96f794;
// music[7917] = 256'ha49a299b239bd09a299563946a975d9714974d962095e595fc939f90098f3c8f;
// music[7918] = 256'h4a96aa9708922496d794ff90439a339d499927989c9309912591d98ecb911895;
// music[7919] = 256'hcb908e93a9987d93309231931891e992c1913e8b5788f48c6991828ec58be48e;
// music[7920] = 256'h2493bf90948c588ec990e6933f943e92e9940590c08782893a8d408f8090b691;
// music[7921] = 256'h518f0d8ace893b8b118cd388d084ee865b871689e388d186568a518a3a8c5d8d;
// music[7922] = 256'h5c8b0b90218baf83f887608db69008934b94ff8dd088628d9b8f3d92f793d393;
// music[7923] = 256'hbb94f8926493a390988fc993b193d394a1920695d0a3f4a93daa7dad9bb088b5;
// music[7924] = 256'hbeb811b8f2b518b456b6e0ba47b9b4b489b4b8b685bca3bf10bcdbba41bb67b9;
// music[7925] = 256'h35b921be71c282c280c37ec03bbbefbc8dc112c207beb4c05ecb73cbdbc443c6;
// music[7926] = 256'h73c6e8c38bc7a8c850c8a8cdecd230d6dfd5fad34cd2e4d405db3ecb93b60cbd;
// music[7927] = 256'hd0c397c1bbc34fc66bca14c9dfbd57ba79c6d2ca47c113c87dda99e188e448e5;
// music[7928] = 256'h98e1aae031e4dde641e36de269ea85ec96e9ddee14f2cdef58f0cfefe0f1abf3;
// music[7929] = 256'h71efdcf11af732fa69ff2600ba024c061d0016ffb3067a06bd05ab0bbc0c9e0e;
// music[7930] = 256'hf911290bd5083d10ae151718aa18a41b721c721a241c7b1c4f1f202341220822;
// music[7931] = 256'hda27ee312a31662fcd364335753478361d348c38fe395d388f3b7f3a1e389939;
// music[7932] = 256'h743bc9392c38b43bf93eb240e1432c430341264578461e4502463a417e401045;
// music[7933] = 256'hb24ae051d2444f36663c143ad332e238ea3f943e9b396b39083dbb3ec73c5b3d;
// music[7934] = 256'hee3f653ec03c513bff3be43ccd36f4338c38e03e013fee37dd3970421442103e;
// music[7935] = 256'h9f410844e53d4c3d54405141cc467f4a31497344f344594b78477944d4487849;
// music[7936] = 256'h304a824820489f4bd04bbd4a92458b49235d9f66bb663468bb664b63f360d966;
// music[7937] = 256'h0e6dd66b0b6c4d682065fc6a0e6ed46ed66d54680969e16d4d6a75618461046a;
// music[7938] = 256'ha36a61657368366aec635c64756684638668476d4e674163e6641564c3639068;
// music[7939] = 256'h4766425e1e6293697b68be657769306d0964be5d446080542f4ab3503351f64b;
// music[7940] = 256'h494b7a4927485749014787418d43234c784b0745eb47f44b8047394379412141;
// music[7941] = 256'hf6448a4633430840dc3ed2403b41ac3f9d43d243623adf380d3fc03eb53b063b;
// music[7942] = 256'h223c163a08382340254100389c3a013d79340f3183360e3ab438433867357532;
// music[7943] = 256'hb73664360e3204363b36ec306f344434f82e8934a1355f2c2c2a4b3257395e33;
// music[7944] = 256'h542d8630d733e435de32972ec52c442be32ef52f712b8124901ea71f7920441f;
// music[7945] = 256'hc21eff202225c520791b651a9c19b419c9167115d115971437124c12c9182812;
// music[7946] = 256'h65064d09af079b076e0d790aa1067000aefc5802d20001f8a2f7b7fe02fdaef6;
// music[7947] = 256'h52f600f327ee36e8d2e252e5b8e78beaa8ea97e7b3e861e3aae153e490deb2e1;
// music[7948] = 256'h64e85de71de625e051dbeae034e798e20fdffde1a9e018e291df4dda3add35d7;
// music[7949] = 256'hf9d40fda55d5b7d562d5e5dad2f5f60467ffacfc58001c03fd004ffd8efdb2ff;
// music[7950] = 256'h16fb00f958ffbefbf4f422fa57ff4cfd11f849f5d2f13beb40ee36f5eaef92e9;
// music[7951] = 256'h06ee78f2aeeff6eeb1ef0eead7e7f5e95de785e6b8e721e709e79de59ce57be5;
// music[7952] = 256'hece149e2f1e3aee262e4a9e460e14be3f6de59cb21c26ec7fbc5ccc4f4c446bf;
// music[7953] = 256'h04c167c307be40bd78bd24bc2bbcb0b71db350b361b4c9b3f1b3e0b6bab540b1;
// music[7954] = 256'hc5b1f4b3e1b307b342afa3ab6bad53b029b5fbb66ead5aab55ad469fea94a296;
// music[7955] = 256'hbc97de986e975e928d8f9a929298c39aca973e96a4983e983b95d591f7909b93;
// music[7956] = 256'h378f918cc691c093fd968c97389384936a91b18d8793499b6999629a9fa224a1;
// music[7957] = 256'haa9d929f659e399f949ddb956f9846a0619eda9c299bf9948398d09900951c9b;
// music[7958] = 256'hca9eb19d679f1e9ba897fe99e39dcaa0399f5e9fcaa3b0a36ca177a47ea862a9;
// music[7959] = 256'hf6a5d49e2c9e16a446a468a1c0a8c2b268b14fad60aac3a6c3a8a0a80fa3f5a1;
// music[7960] = 256'h18a61ea956a98daaeba9b4a7bbaad5ad2cad34af45b272ae45adb0b68eba33b6;
// music[7961] = 256'h52b68eb9d9b957b986ba1cbad6ba34bc7eb97abac1bdc6bcc2bb19bee2c1e3c1;
// music[7962] = 256'h9bc19dc384c5f4cd73d8b2dc32dfbae13de273e184e212e545e5f7e44de756e9;
// music[7963] = 256'h96e715e6cee706e958e7e9e681ea8fedd9eefcef5bf0ebeed1ebe9ea99e922eb;
// music[7964] = 256'h56f1b9f0e7ed06ee99f324fb2bf6dcf3fbf56df570fcdbfa36fa9a026a00d201;
// music[7965] = 256'ha9ff92f694fd470176ff36061400eded38e755e9f2edb6f22eefd1ea7eeb4eeb;
// music[7966] = 256'h95edfaeea3ece5ec85f0f6f022ee95f0a7f301f5c6f7a2f6c4f638f6a0f249f7;
// music[7967] = 256'h5a00920247ff93fb3af8c9fe32075cffc3fe22050f015d02a102e2022a081105;
// music[7968] = 256'h83066e092d04f30311067b0aa00f610cdd09610bb70b1b0d190d030eff10570f;
// music[7969] = 256'h48109514a0137a1334145f146918261cee1b7e1a7d1bd41ff52385221e232d2c;
// music[7970] = 256'hc12de02be02f0a2e5c2b2a2ccc2b042b3e296a2a802e5232a430a12f35351333;
// music[7971] = 256'h7436da44fa48e64ab34b774ae74cf849054a2c4c214a8f4d654f234c1f4bdf4c;
// music[7972] = 256'heb4f0e5183528554a752414e014da34f7650754eba4d47506352b0523d547750;
// music[7973] = 256'h35490649844a0549e848384a704a474ed751cf4cd04e88544b509b5274555a52;
// music[7974] = 256'hfb52494fbb4d07518b509d50244fcb4dbc4e6350da52d95277525c507e4dd54a;
// music[7975] = 256'hc04a8859b768896b3f6c5c679860b860bc617a5f7a5f5e63886342601c5e6561;
// music[7976] = 256'h9467c964aa621c66dd63a9632066095d474e0d48d946cf4453454948684c344c;
// music[7977] = 256'h2d466b4277429644754587438c416540cc4279454346b946f7447543603f5e3b;
// music[7978] = 256'h65409b41ed3d2e4197388825102213222f1f531f671cc7217524941a721b9d1e;
// music[7979] = 256'ha21aec1a401e1b20d61cca1995186d16d71698157e1234129a16fa1a1e195f1a;
// music[7980] = 256'hd61ca9178312c413fd17fd188316e411ca0f691304123b0ef20e2f0fc4104d13;
// music[7981] = 256'hf4121110d80ed312bf12440c680da013ef0e0209cd0dd2101a0f0d0c49068206;
// music[7982] = 256'hcb0c3d0ea60ce80e8010f30e100efc0c360cb50af90acb0e860d840b450fc413;
// music[7983] = 256'h9d13220cf00acf11990fc70a6c0e1f11b60f1313dd156111a70f7d0f6d0d4d0e;
// music[7984] = 256'hdb0f9a112c114c0e820c4709fb073908db06f7077208d4064d08a4092d060f04;
// music[7985] = 256'h2d052005d7078e07b8fe73fb3ffffa00bfff39fda0fc2dfd47fc37f91bf719fa;
// music[7986] = 256'h39fb26f776f46ff44df555f601f625f3d8f0aff12df15bee26ef7ff4c3f636f3;
// music[7987] = 256'hd1f06cf181f296f34cf2e1ed8dec24f1e2f258f0aaee29edcdedafeb1bec74fd;
// music[7988] = 256'h140c0f0b480aef0a6807b600abfd1c00ac00ff015a0334020e0241fffffd6801;
// music[7989] = 256'h990110ff98fee800c40128012b01e4fdc7f920f9f0f96ef8f1f503f831fa62f9;
// music[7990] = 256'ha0f90ffc3afde2f848f687f631f7a3fbc0f7b6f0fdf48df7b2f344f202f542f2;
// music[7991] = 256'hfeee0bf69aecaad7f3d727dc14dc94dcded713d7f3d601d573d600d5cad331d6;
// music[7992] = 256'he4d964dbf9d785d737d9a0d753d54fd3f6d30ed21dd0fedca4eab2ec57ed77ea;
// music[7993] = 256'h4ce862e99fe5bae596e6fee3e4e70ee9c2e40ce36ee297e2b6e1d9e20fe54fe5;
// music[7994] = 256'h6ce73be5f9e122e476e44be3c7e2f6e49be7d6e679e653e24fdea6e1cae434e3;
// music[7995] = 256'h69de51de56e1c7de6ddfd5e6b2eab3e77de8cfeb74e8e8e8cfe9f2e88cefb8ee;
// music[7996] = 256'hd4eb1eeeb0ea3dedf5f0b3eecdf102f1c8eb27eb2aec50f15cf558f1bded16ed;
// music[7997] = 256'h88ed4def55ecf8e965ed1bec9ae905ed41efe8efaff040ee9aeb9eecffeb21e9;
// music[7998] = 256'h83ec5ded96e173dc7fe0d8da9fd733dc09da92d80ad9a8d64ad7c0d7fbd790d8;
// music[7999] = 256'h55d58bd4d2d7ddd6ffd488d8f8d897d8f1dac0d580d273d469d280d6d1db45d9;
// music[8000] = 256'h6fd85ed8ead6ced94edd58dcb4dadbdaefd9cbdabdda9bd29dd802f4ccfd95f6;
// music[8001] = 256'h2ff641f548f3f1ef3feeb8f435f8dbf67bf130ef31f393f17ef107f442f4a8f4;
// music[8002] = 256'h78f227f21cf0d3ef55f479f2d7efbaed8aec01edbeeba6ef47f1f6ee53efc8ef;
// music[8003] = 256'h2bf287f078eb60ea86efe5f148eb90ec9cf032ef70f049ed10ec2eeb51eab5ee;
// music[8004] = 256'h2ce1c3ce04d192d8e8d6cdcdf0cecdd409d0cbcf96d291ce42cbbfcd82d1a8cf;
// music[8005] = 256'h71d2c3d78cd29fcf6fd1b8d3c9d74fd303ce33cf50cefbcda3cd39cd5bce83cd;
// music[8006] = 256'hd2d00ed5dbd2bbd0eecf4ed288d775d510d39ad616d5e8d29cd44fd178ce7bd1;
// music[8007] = 256'hb1d43ad529d575d787d5a5cef4ce54d449d6edd634d7ebd3c2cf1bcf8ccff5d0;
// music[8008] = 256'h4ad3a1ce55cbdad311d5a1ce59d28fd5afd6ced845d496d220d3e9d164d579d7;
// music[8009] = 256'h1bd8ced811d5a1d3bed8c4da4ed869db39de28dbded9c3d804d8ebd901dab3d8;
// music[8010] = 256'hdad871daa2db25da7fd73ed8abd981dac4dd28dddcd90cd809d738db37e0dae2;
// music[8011] = 256'h0ce2b9de64df77dc9bd7a8db26e02eddebd846d951d982dbd0df83de97de26de;
// music[8012] = 256'h25dc7be084e032dceedb63dce5dc0edd40db21dceae13ee4eae2bde417e6a9e8;
// music[8013] = 256'he9ecc0eb1de81ae8b1eba2eee4ed17ee4feeffeacaf30507ae0a87091d0fe60d;
// music[8014] = 256'h690b850b760b7d0bb809c010d91ea4245523622188202223432591225f229a25;
// music[8015] = 256'h61279a28ec27af26512596258627da26662ae42c9a29fe29ad2af72a7b2a322a;
// music[8016] = 256'h022e7e2c8f2a512b5a299b2b452ed52eac3054305a2e162ec2339231341f9a15;
// music[8017] = 256'h6519ff1aab1bdd1ce91abd177f18011b571bc91c7a1ea01d231c071b031af81e;
// music[8018] = 256'h2d24141e551e72233a1f4f22d2214f1dbe22561eec1d6125a122d123ef22ec1f;
// music[8019] = 256'hdf23d322112200237921da22de238522f823cc2596243224831cb0106412e513;
// music[8020] = 256'hea101c151f175a1589168a189419ea17fa122e102b1373176c1ad41ce91f261f;
// music[8021] = 256'he41bad1d271f7b205921f11e7322bb2440222e222f227f21691f9a1f88211d24;
// music[8022] = 256'h892c66300a2efe2dd82cb82aa52b012df82bf62a6a2be62e4c31b72c2a2a4e2b;
// music[8023] = 256'h3b2d90310a322730842e482c152f3933f62ed929562eb0316630cd30f12e2b2e;
// music[8024] = 256'h8030da30b12dd6290b2a6c2b492b9a29612a8d2f412e492a362ce32d2e2e092f;
// music[8025] = 256'h1d2edd2a3b28782728285c29712851289b29e52811268b26932b552c592ab929;
// music[8026] = 256'h8429812c4b2de42b182de22fb22eea2a7536f846e046a3453549c34715440d43;
// music[8027] = 256'hf443da43ef43b144bc434a44a9470448ce45e145474432409e40d3463d498f47;
// music[8028] = 256'he548e5466545544655429545344a7448874a4a498247c648fa459745b8437940;
// music[8029] = 256'h6444f0434a3f734190433244ef447143bf40933c5b405440df2dce26d92cfb2a;
// music[8030] = 256'h2228be26aa27bc281926f923cd22b42270244d297e29c2243b258c2531278227;
// music[8031] = 256'h34244f25e32382234825a521551fd81f49236d2383211223ce1fda1eb220f41e;
// music[8032] = 256'hf2201521561f3e1f5d1c8b1b221e4d1f4e1fbf1e3a1d7f1c401d1e1cec19f519;
// music[8033] = 256'hb919fd16a313f01025141519fe156c15c7177f14931511170414ff14cf155014;
// music[8034] = 256'hf2142415d01458166515bc12f914e716351631169614c115ff193d1a5f18cb17;
// music[8035] = 256'h4117d5154d16b418e9189318c417be13b40e420da5133816ff10e31241124711;
// music[8036] = 256'h3a1e57248f227b21fa1d2120c51f641d881e5a1d2e20a71e1f18fb178f18ce18;
// music[8037] = 256'h9516941367134612a80f6e0cae0f4d12a40ea5106a10420d8d0ce0081109330a;
// music[8038] = 256'h67081409910717044a020005aa083806eb06bb087e026c01950373019f049605;
// music[8039] = 256'h0602930172fddefddb02abffc5051d17a81bb315eb12b313ac139d122911870e;
// music[8040] = 256'ha00d600d8c0dcc0e5b0b7b0ba30e8a0854072d0b2907c5037303de06d9079702;
// music[8041] = 256'hf40488075e03c1ff2ffe1502b7febbf0e2e9f3e8cee7bce65ce58ee59fe695e8;
// music[8042] = 256'h68ea5ee7cfe1c5e0c0e1a7e2fbe37de395e336ddefcf54c917c897c910ca07c7;
// music[8043] = 256'h54c745c745c738c8aec656c554c317c46cc5e0c3b2c559c497c0eac0dec007c4;
// music[8044] = 256'hfec52ac1edc1b7c385c095c295c2ccbedfbf9cbe17be7bc052c0debf9bbd07bd;
// music[8045] = 256'h14be20bca3bb74bc85be31bf16bdb8bc3fbd66be11bd2bbb4bbc69bb37bb7dba;
// music[8046] = 256'h1ab9c4bc00beb1b98fb680b7d3b951bb96bba2b98cb9d1b912b844b989ba2cbb;
// music[8047] = 256'habbb5abab0bad8b94eb709b893bbdebebfbd50bd55c0dfbec0bd77bf15be23bf;
// music[8048] = 256'hbec1b8c2dbc39fc0cdbea0c1c4bfb4bdcac0e2c1a7c09ac1c1c1cdc1f3c2d9c0;
// music[8049] = 256'h22c021c1ddbea6bef4c2fac6f2c3d1c097c325c2b5c0b2c2a8c301c493be0cbc;
// music[8050] = 256'h16be78bbbebc4fc1cbc327c563c3b6c21ec294c052c14ac105c1d5bf66bd11bf;
// music[8051] = 256'h66bf89bd54bfa0bf1abfa7beacbd26c13bc166bfd9c21fc53cc66cc558c437c5;
// music[8052] = 256'h49c82fd13bd054cc49db36e6ede23ae1a3e071e0f0e128e5c7e83fe990ea90ed;
// music[8053] = 256'h13ef9ff0f4f04ff332f88bf74cf85ffad5f50df526f533f2a3f4eff55af6f9f7;
// music[8054] = 256'hc0f4f1f262f35bf15ef0fff0c7f08fee58eef1f01dee89eb37ee94ec43ebd2ea;
// music[8055] = 256'h17e71ae74ee7e5e7bbe812e85aea4ddff5cd6bcd03cf58ccc4ccb0cb48caeacb;
// music[8056] = 256'hc3cdbecd4fce63ce90cee6cf0ad0f7d0efd16fd2ead211d1fed052d4ecd55ad3;
// music[8057] = 256'hfdd314d74dd6b7d7e4d81cd801d92ad93cda95d9d1df1fedbfef60eeddefc7f2;
// music[8058] = 256'h81f42bf2f7f48af689f43ef628f59df56af8a0f880f9c7f936fae1fa9ef9faf7;
// music[8059] = 256'h33f81afaf5f9d8f91afbd8fbcafd14fe22fd1d00e4013b00c8019204ca046f06;
// music[8060] = 256'h9707e405500784091909f20c9a0f780c760d0c1095103f12da1219138b12f512;
// music[8061] = 256'h9e15011723180a187b17dc1793171b19fb191319c419671b8e1a9518581a5a1c;
// music[8062] = 256'h8c1d751f7c1dff1a5a1b5c1c7a1dd11f7b20621e491fe81e411e70216020bb21;
// music[8063] = 256'h9b20041222086009730bc80b920c7c0c7709360b8e0e230d0b0efb0e4b0dee0f;
// music[8064] = 256'h9213c1111411c311770f791088118d10ea11ed1110131c146b13b813da14fc17;
// music[8065] = 256'h5215e1163328e72f752cf32e3530f42ee52f0030e32fde322f3551344134e333;
// music[8066] = 256'h4b336d333e33f0323c3176329c34f533d735243570325534c934cb33f133de32;
// music[8067] = 256'hd6309f312a350b349632783465336d333d331f31bf31223181311532fb2f8130;
// music[8068] = 256'h9f3089302131ed312b33e82775182616cf16781796198d1752171b196017d016;
// music[8069] = 256'h921785174519bc1858179e18c2170d18cf183b17fd16c9168418c118b3161519;
// music[8070] = 256'h78190919c11be31b0a18f4124a13a315a2157c19751db41d661c111c341cc61a;
// music[8071] = 256'hdf19aa1669135214ac13c313e014ee1257126512b10f1e10b213801284114414;
// music[8072] = 256'h5914c61469153114c416221b8f1b1c1b1f1d201c1f1aa11a3119e41b9c202120;
// music[8073] = 256'h912135240e274f2a392aa52a792b202cd62e603041306930f130f13095308630;
// music[8074] = 256'h2c31c430452fd8308331762f9b2f392e072d852e262d212ba42b0e2cba2a4a29;
// music[8075] = 256'h2528c425fe24d32511266426c225e6244823b620fc20e021cf20381f5f1e301f;
// music[8076] = 256'h321dc118fd171318531658141c14c215b914241228122513c311dc0e1a0fa90f;
// music[8077] = 256'hf30d6b0d6d0d120c140ad009960932097e0ace0819075606130682088504b606;
// music[8078] = 256'hda166a1bd5160c18f019b81944184b188418a716cc14f2128613e31493121a12;
// music[8079] = 256'h48131c11350f800cd70ddd1aaf220921d422bf2235215822b520161f051f3f1e;
// music[8080] = 256'h3c1d731c691cec1a3519311a5c1ae618a81708170c175615d8135b1481156e17;
// music[8081] = 256'he8152d16ce15030699f8f4f8fdf8aafa50fb44f917fa9cf910f946f91af895f7;
// music[8082] = 256'h91f8d3f95bf87cf722f93bfaa3f95ff735f711f9c4f810f81ffa58fb0ff92af9;
// music[8083] = 256'h45fadaf9d4fa48fabef803f830f84bf9a0f8a5f8fcf974f98ef672f574f8ddf8;
// music[8084] = 256'hf5f740f9fdf8faf7bff808fa1ff8f3f768f9a4f697f8b8f4bce5c6e2e1e401e2;
// music[8085] = 256'h42e384e4cfe4d0e4aee3cde428e595e4e7e497e556e7c8e63ee6ace84de940eb;
// music[8086] = 256'hfdee0bee5eec96ece7eb30eba4ea52ea97eb62edb8edc7ed0fee1eed7fec3bed;
// music[8087] = 256'h2eef97f09eef8bed53ee37f3f4f28eefdcf223f3a1f0ccf155f048ef97efc4ee;
// music[8088] = 256'hb6efa7ef89ee39ee03ee39ee07ee97edfeed1fef4fef87ed7aed56f0ccf04ef0;
// music[8089] = 256'h2bf1afee66ec78eb8fe957eb38ec8feaebea2eeb16ecc5ec1dec32ecbdeb6eea;
// music[8090] = 256'h15eab4eb38ecc3eabbe992e94be94be761e62be839ea56e8aee477ef70005b03;
// music[8091] = 256'hf301cf02d001d6019e0296021602dc018d0149027f03f20255023a02cf027f03;
// music[8092] = 256'h0e02ad002b022b042003ce02520350022b03f7021c02a402cf009400b901ee00;
// music[8093] = 256'h2501cb019701e10060009e01da027b02ec01fe01670201026701fe0183019c02;
// music[8094] = 256'h0800dbf0d5e558e6ede682e76be751e783e8dbe8fae81de818e807e819e875e9;
// music[8095] = 256'h14e971e91fe9e8e78be8d6e7b7e745e83ce804e83fe7c9e73ee868e8b3e885e8;
// music[8096] = 256'h37e97ae9e2e87ce7e6e650e795e7e6e70ce74ae73be8d6e827ea5ae900eac3ea;
// music[8097] = 256'h7ce95dea2ceacee9bbea3eea51eae3e92ce97ce99ce986e9d0e98beaebeacfea;
// music[8098] = 256'h7aea3eea60ea67ea2feabde954ea2beb57eb9aebfeeb08eccbeba6ee71f2e1f1;
// music[8099] = 256'h87f07cf086f028f09def40ef8fee20ef7eef58ee33ee99ee56eeacee8df06ff1;
// music[8100] = 256'h97f17ef158f14ff4e4f5b9f458f409f41af442f3e5f252f23ff2e2f2f4ef2cf7;
// music[8101] = 256'h61053307cd057e07be08360917087008450824085a080a07060725070107e007;
// music[8102] = 256'h8507fc03da00fe019102c102fc03fa0368040b04e5021d033a033c0368033d03;
// music[8103] = 256'h1d0300030f010a009600b9ff1affdefd73fee8fea7fdb309b71857196b183719;
// music[8104] = 256'h99183c197a18351897189318ac19a0190e196619c8180418d41769179b17fb17;
// music[8105] = 256'he217d517cf17b817211715178b177617bc1760171d16c614f113ef13e6125512;
// music[8106] = 256'h9c12651295129311d112dd12b6074cfefefe0efe24fdd6fca0faadfdfef8f3e7;
// music[8107] = 256'h55e100e37ce236e34de397e306e496e316e465e32fe395e32ee339e3fae2c2e2;
// music[8108] = 256'h56e205e23de20de22fe200e2c7e17de152e1f3e1a1e162e119e272e200e2b6e1;
// music[8109] = 256'hfde24be3a5e2c3e226e2c6e1f2e1eae1b3e19ae141e23fe294e1f5e0c9e056e1;
// music[8110] = 256'h46e122e158e11de22de3aee222e26be284e2a3e252e227e22ee20ce254e26ee2;
// music[8111] = 256'h79e29ce278e277e25ee276e29ee239e28be259e386e35be4abe57ae654e78be7;
// music[8112] = 256'h00e7c2e642e690e51ae55ee446e48ee4c3e389e3b0e35fe3e3e413e79ae8ece9;
// music[8113] = 256'h55e952e852e802e8dde7d3e79fe751e7e0e6c0e685e6b2e630e798e7a0e8fee8;
// music[8114] = 256'h02e99de95de9f0e8f5e80be904e9cde76ee704e9a0e943ea2bec91eb9de776e5;
// music[8115] = 256'h22e798e84ae9bdea20ec58ed21ed4bec42eb17e9dfe889e970e923e95fe80ce9;
// music[8116] = 256'hdee79ae469e308e4cee5eae5dbe6b4e6e3e6b4f590034a02f8015803ae06a60c;
// music[8117] = 256'h990bb809710ae6086e0803094209af0a460c3b0d8e0e4b10f2117d1303154716;
// music[8118] = 256'hc1177419681a221b961b5b1b641b471b791bd91b981b5a1b8f1aba195f197918;
// music[8119] = 256'h54189518e0177c17a9167f15c715af1457146a148b128914c10d1cfc6bf7f5f8;
// music[8120] = 256'hc7f6e8f67af6b2f6cef617f66df6baf5c1f5eaf4f0f3e4f3d2f201f34cf38ef3;
// music[8121] = 256'hdcf3eef22af25bf15ef161f11af131f1dbf09cf116f2aaf1eff11ef223f2d4f2;
// music[8122] = 256'h83f34af4c3f6a3f75df72cf84cf708f80bf7bff859062e0e8e0c4d0d750d550e;
// music[8123] = 256'h090f260edd0e120f4a0f6910931073106710d90fa20ffe0fef0fe11087110b11;
// music[8124] = 256'hf8106d100d103410d80fb90f71103c1163119d1123123f14f714cf1212141616;
// music[8125] = 256'hd015a51651169015a515f114bd14351501157f153a18bf1ad51bfb1b6c1b5c1b;
// music[8126] = 256'hc31af71ad71bbb1b111cb41b951bbd1b5b1b581cfa1c391d4d1d3f1dd41dc11d;
// music[8127] = 256'hc11d011dcb1ca91daf1de71e3a1f7a1ec01e1a1ef01cf21bd71c811c951a381b;
// music[8128] = 256'hcf1430094006ec055104dd04a1033d03cc043204f304a60556044e04a3037f02;
// music[8129] = 256'h7b020204f4048a03d004d3035005c714d81e261d311ead1e671e931f7a1f1b20;
// music[8130] = 256'h772070206621d921ce2163216921df21c121f6218021ef20c1222a243324b424;
// music[8131] = 256'h8624e12396233f230b23202381234923d0225e23b023c822fa216a2120219120;
// music[8132] = 256'h3d1fb91ee71d1c1ea61fd71ead1f2c1f051e90206416db06aa05e0065f069207;
// music[8133] = 256'ha207c208aa099c095b092509de08d107fb072e086e084b09de08c408c3084508;
// music[8134] = 256'h8008c8089508470880086c080f084c083d080408e2079f07c3073d08e6084b0a;
// music[8135] = 256'h300d620ebe0729015505b5099b0a110fe6104a11f7128f118610240f860c3c0b;
// music[8136] = 256'h8a095d0866078805b8038b032a0476033e047805ff05c7077408e5092b0b560a;
// music[8137] = 256'h150bf70bf50e2715ae1627154216f316ac167118921ab41bc91cdc1d3820c723;
// music[8138] = 256'hb825cd26c428aa298a2a212d4b2ed52d3f2e6930f13151315131e13029308730;
// music[8139] = 256'h622f822e682e5a2ff630602f262eda2de32b852a87290329b8284428f9277a27;
// music[8140] = 256'ha4274227c62643264925ca24c523ca223021f51fac1fed1daa1d311cf9180118;
// music[8141] = 256'h69162a153f1387113513be11cf0e0b0dac094b08a308c50729066e049a030504;
// music[8142] = 256'h2a037002b903020159044e14b01a9717ec17a3165415c614e3121412b710540f;
// music[8143] = 256'h630e130da50b290ac009ef08fc0660050f049c03fb02a1011f014b007dff88ff;
// music[8144] = 256'h96fe8aff35ff2cfc3204cb0fbb0f520e1c0e490d4f0f570e940c810c050bfe0a;
// music[8145] = 256'h6b0a5109b008c806180764062906a3064df911eb25ebc2ea98e992ea3ce9b9e9;
// music[8146] = 256'h08e99ee7dee7c5e68fe69ce669e66ee694e537e59ae466e486e4e0e379e3e4e2;
// music[8147] = 256'h66e2dbe18ee19de14ae105e144e0a1dfdade61de1edf2bdf88dff5dff5df81e0;
// music[8148] = 256'hafe00ce137e14be187e152e1b2e19ee17fe160e13fe1a5e135e12be187e1e2e1;
// music[8149] = 256'h5be286e22de378e2cce242e38ce2bbe3d6e174e179e0e7d3e9cb3fcde5cc11cd;
// music[8150] = 256'hbbcb97cae9cbafcb1bcc66cc16cca0cc47cc64cd5acf16cfe8cec3cee7cd9ecf;
// music[8151] = 256'h8ad2b9d2c2d152d16bd038d0f2d14cd3e1d270d26fd20ad29ed195d1dbd13cd2;
// music[8152] = 256'h4fd284d21bd37bd305d434d4dad310d4f9d3b6d4c8d613d794d694d604d691d6;
// music[8153] = 256'h8fd7bed62cd65bd6d7d59dd57bd5f8d4b5d4ced4e3d4b7d427d537d426d257d2;
// music[8154] = 256'h8cd243d3c8d3a5d043cf59d116d278d210d4d8d39bd236d324d3bed32bd41fd4;
// music[8155] = 256'he6d520d49fda92eb69ef2bedc3ee5eed4feddaeda9ed99eeb7eef5eecaeed5ee;
// music[8156] = 256'hd6ee45ee97ee72ee5fee16efb4ef55f0d7f03bf130f16ef1bcf1e9f1c2f2d6f2;
// music[8157] = 256'hbef24df3a5f367f4f5f4f2f4aaf429f4dff3d7f393f4ddf49bf432f5edf483f5;
// music[8158] = 256'h8bf558f3baf3d9f3f7f4daf397e5a9db3ade6bdef3deafe07ce011e108e197e1;
// music[8159] = 256'h5be287e2dde2a1e2c7e214e347e369e3b8e332e418e414e483e36ae3ece3cde3;
// music[8160] = 256'h2de401e4c8e3eae3cde3dbe338e378e313e438e47ce5e7e508e606e795e71ee8;
// music[8161] = 256'hd3e82fe990e9f3e9f3e997ea1debe3eae7ebbfec3eed36ee94eec5eef8ee69ef;
// music[8162] = 256'hb8ef1bf0def0c3f031f1b3f199f1f2f1d6f196f1fff150f204f22df20bf35bf3;
// music[8163] = 256'he3f3dff381f3fcf325f440f4aef4bff4e9f4c2f6baf826f93efa63f912f8eef9;
// music[8164] = 256'h88fab6f974f979fa14fc83fbeefac4fa9afaabfa56fa98faa7fa20fbcffbeefb;
// music[8165] = 256'h89fc02fdd8fd7ffefafe23ff0fff0b0079ff97ffeeffe6fe45000dff83024411;
// music[8166] = 256'h2818ba15fd16e0180a1978193019d318cc181b199a192e195919a31831155b14;
// music[8167] = 256'h8d153016f316c9154d15ee169b1642151016f6169b164b17da167217ee172615;
// music[8168] = 256'h921e622ef82f672e592f152ea32e752ed22d582e292e702e382ed82da72df82c;
// music[8169] = 256'hf22cb52cc02c2c2dec2c3b2d8d2da92d0c2e002ee22dc12d6f2d532db62df22d;
// music[8170] = 256'hf12d982eb82e332edd2d952d962d542d272d242d652d7c2d622c712c832cf02c;
// music[8171] = 256'h1f2e2f2d732e272bb21bad0b370166fee2ffc6fd9cfc69fd94fd28fe01fef0fd;
// music[8172] = 256'hb9fd9cfde3fd9efde4fdd7fd64fd1cfd84fc1efceefb00fc14fc40fc82fc59fc;
// music[8173] = 256'h4afcebfb4afb36fba9fbd8fb8afb9dfbbffb3cfc10fd19fd60fde3fd36feedfe;
// music[8174] = 256'h30ffeafe65ffe9ffd9ff07018002fd02ce036f032b020002da012a013e00cfff;
// music[8175] = 256'he2ffeaff3f005e00a2001701bd00030075ff43ff81ff82ff4bff98ffbbff9aff;
// music[8176] = 256'heaffbbffaaffb2ffb1ff2500550043026c03cf029b045704aa025202c5000403;
// music[8177] = 256'h0a06e7045204c203230375030c03bd027c021902d601a4018b01fc01a8027102;
// music[8178] = 256'h72029f02990267036303c602360387036003980395033e037903e303f503d003;
// music[8179] = 256'h7b032003e702e5027a029a020603c50220032a03a902f4ff5afa45f9d1fb1efc;
// music[8180] = 256'h8cfd8f019f02b3ffdbfed7ffaaff44ff65febbfda3fc9afcaafb9cfad706fb13;
// music[8181] = 256'he812f411ea12781250137112661214136013c4136912d712df17e51bc1197717;
// music[8182] = 256'hb217f7150116c9165c16e5173c19071b011d0b1e0c205621b5223824d324df25;
// music[8183] = 256'h782611276e277327af270e27c1266726da257025d8247525702419239222d120;
// music[8184] = 256'h7f222e1c8d0a5204f60553048f04770339029e0222012500a4ffb1fe05fe93fd;
// music[8185] = 256'hfcfc8bfb98faf7f964f9b9f885f72cf7c7f640f651f6ddf5d6f5adf677f6a7f4;
// music[8186] = 256'hacf36ff341f2c2f19cf143f178f162f126f170f102f224f26df29df24bf2cef2;
// music[8187] = 256'hecf204f3fff274f2ccf222f268f2b9f170f0bdfa9a06a60768084309d707be07;
// music[8188] = 256'h830753081f09d3082409ab080d089b07120767074807ac060b064c05c6043504;
// music[8189] = 256'hd1031b034603100555052104a4035003680209028c02ac02cc02e80284030605;
// music[8190] = 256'h8a04d0033b043e03af02a00225025c021c02ba01bc01dc01140260025903b303;
// music[8191] = 256'hb0030904a503c403f80390039e033f03b9028402490235023802470258019200;
// music[8192] = 256'h0d01eb00ba00ea001f01b70078fe0ffd7afdb7fd66fd88fd2afe2bfd41fcbff6;
// music[8193] = 256'h6fe824e117e2eddfccdf6ae02ae025e145e09ce179e090e020efccf9f8f77bf8;
// music[8194] = 256'hfef8fbf710f8f0f6a2f685f650f6a8f68bf638f774f754f7e9f7b4f73cf7e6f6;
// music[8195] = 256'h03f703f7a8f60bf750f6c1f518f695f5caf5a6f55af5e4f516f69ff7c8f887f7;
// music[8196] = 256'h40f646f61ef661f5a9f531f58df5bbf669f513f5b5f406f4a2f39ff263f447eb;
// music[8197] = 256'h13da6cd743d982d7d4d7dad605d77ed7e5d670d77dd791d76fd7ecd682d6d1d6;
// music[8198] = 256'h2fd815d840d7a9d637d6abd66ad6ffd5bfd66ad7a0d7f5d7cdd786d7b7d7a2d7;
// music[8199] = 256'h0bd87bd899d8fcd860d851d8b1d8bdd847d937d9c7d924da2eda39dc1fdf3bdf;
// music[8200] = 256'h37d788d125d7afda5adc5ae1ece2eae3cde428e35ae229e176df29de4adc09db;
// music[8201] = 256'hfbd96ad9f0d8e9d695d6f2d7acd857da48dbb6db64dd93de29e02ce166e0bce1;
// music[8202] = 256'h12e770ec3fed83ec00edb0ec73ec9eed82f04ff3d5f5b9f9dffbd9fd6e01ee02;
// music[8203] = 256'h3b047706ed07ea08e1092c0b090cd00c180efd0ea70fe10fe70f8310c410960f;
// music[8204] = 256'h880f1f120813d711a211a6106c0f290f110e810d570da10c290da60dca0d990e;
// music[8205] = 256'h340f570fe90d5d0cfe0cfc0d100ec60db90d290d2b0c850ad3085d09ed078004;
// music[8206] = 256'hc203ea037d045403350232024700a400f4fd64ff2c104c1835154e166015ac14;
// music[8207] = 256'h7815c214ca152e169115671566157b1573155e1517145813f612ee118511d310;
// music[8208] = 256'h0a10e70f1a10a80f8d0ef80de00cb00c070d9e0c900c1a0c200ca90b4b0b740b;
// music[8209] = 256'h7b0ace0bc90b0e10231d9e20ea1e5920b61e16212d21a31f352255166b076107;
// music[8210] = 256'h0f0825078807b306e206c506c206f906ba062e07a40622066f0637069306a406;
// music[8211] = 256'h12061206c505a905510658064006d906a806580605077607f5076108fa07c707;
// music[8212] = 256'h00084808b20836095c098c095a0aa00ad80a500ba10b920c4d0d780d200ddc0c;
// music[8213] = 256'h910df90daf0eff0edf0eb60fac0f1010af10d2101512e011c911771264120c13;
// music[8214] = 256'h2413bc133014dd145f16cd15f316b915df132e16be0c380202055f0585046004;
// music[8215] = 256'h8401010247026203ff0564051b052405c9041c0507054307bd0a0a0bc309b209;
// music[8216] = 256'h5d09840860083808890820093409410937098309d809210aaa0a910a8f0aba0a;
// music[8217] = 256'haf0ab40acc0a460b920bc90c6f0e180ed70da80d030d480db00cb10cd10ca20a;
// music[8218] = 256'h8d0ad80b970b9f0bda0b970d1e0e3c0be00a650b5b0ac70abe0ab50aff0a9208;
// music[8219] = 256'h690516058806e10569060808d404450afb1a7a20ec1d0a1f671e2b1ed41eb91d;
// music[8220] = 256'h2e1e391ec71d911e8e1e4e1e341e2a1efb1d721d1f1d721c7a1cbb1c5c1c921c;
// music[8221] = 256'hf91bf71af61ac41a991a9e1af81995190d1ac4199c190d1a9c1989193e19ed18;
// music[8222] = 256'h4519b718c4186718f517fd17c3166f17b216d416971776091efb8dfc1bfd98fb;
// music[8223] = 256'hb2fcb8fbcefba7fca4fbe9fad9fa98fa6bfa3bfaf9f985fa10fa55f86ef75ef7;
// music[8224] = 256'hcef7d2f7dcf7e3f775f7e5f7d0f7cff756f8b9f7bff7c0f73df74df71af7c7f6;
// music[8225] = 256'h49f62ff611f6b2f5f7f539f5aef474f4a8f32df407f481f3eef362f38bf317f4;
// music[8226] = 256'h88f36df3aff3baf3b9f3a2f334f3eaf250f377f325f3e9f2dcf29ff25bf258f2;
// music[8227] = 256'h44f2dff24bf31cf345f38ef23cf2c8f2dcf230f470f4d5f2a0f244f2d6f15ff3;
// music[8228] = 256'ha7f400f46ff38ef3baf26cf23df2f9f070f1f9f1a7f2c1f5a7f638f5b7f43bf4;
// music[8229] = 256'he9f34cf358f2d0f12cf1bef08df086f099f039f0b9ef99efbfefaaefa1ef26ef;
// music[8230] = 256'ha5eea7efceef3bef80ef44ef89efdeefa9f023f2c7f1adf157ef8bee4ef9ab02;
// music[8231] = 256'h4f02cb01a400b8ff8c0137020f02e301ac012c017c00da00ba001c001cfe68fb;
// music[8232] = 256'hb1fa4ff942fa7cfbeaf8d5013d1164136d113b12ac11fc117711a4104f111f11;
// music[8233] = 256'h2511b41132118c104410b40fdb0f2a108b0fe70f4310a60fc60f920f450f650f;
// music[8234] = 256'h9d0ea60ddc0d430ed70d050ee80d430de70db00d6f0de30d620d920d5c0d160d;
// music[8235] = 256'h150d1c0c570c0b0cbf0c2b0e820c780efc0b2cfc43f33af52ff426f3b6f216f1;
// music[8236] = 256'h7df21df2c9f080f362effce3b3dfe2e05ce05de088e0dade59ded0de08deb0de;
// music[8237] = 256'h67df0cdf22e0e6df75df13e036df91dfb7dfdcde5edf06df64df35e0c9df70e0;
// music[8238] = 256'h7ae027e074e0d9df00e037e0cddf10e0b3df73df41e013e01ae015e13fe1a4e2;
// music[8239] = 256'ha6e337e2abe2f1e206e2b1e219e20ee22fe3e5e221e330e3fce20ae325e37ae3;
// music[8240] = 256'h13e3d2e3b1e311e300e548e563e6d5e75ee598e577e7e3e7aee82de808e89ae7;
// music[8241] = 256'h28e634e679e690e670e65ee6a9e6fbe67de876e93be913eae0eb46ec09ebc5ea;
// music[8242] = 256'h69eab0e9f1e9f1e873e8bfe840e883e84ce80fe861e831e899e8ffe86ee999e9;
// music[8243] = 256'h56e9cae9cde941ea0aebe7ea50ebb1eb9debc9ea5de9ffe9d5ea5de9a9e80fea;
// music[8244] = 256'ha0ea60eafaea6aeb03eb50ea0dea5eebc7ed22ecbae6dde6b1e849e8c4eb9eec;
// music[8245] = 256'ha6eb5cec9bebc3f63b057904c4020004630209027001a800bbff1bff2f0001ff;
// music[8246] = 256'h5afdeafda0fe5bff6c001d019601f9012d019c02dc08610c910af6082d081207;
// music[8247] = 256'h4207e8073c08460a5e0c330eb210ea113b144e16e516ef180319a4195b1bb61a;
// music[8248] = 256'h531cde1c6a1cbb1d421c391d9819f00a9c04a306f10337029d022d0117013601;
// music[8249] = 256'hd7ff1d00e3ff90fedafed5fdc2fce3fc1efb1ffab7f964f8abf85ff863f7f6f7;
// music[8250] = 256'hedf741f769f74ef7b3f639f6aff54cf567f546f530f5c1f5b3f5f7f4d7f477f4;
// music[8251] = 256'h0af42ef4c7f3ccf397f3b1f22ef38cf319f40cf50bf5eef5e8f50bf60cf872f8;
// music[8252] = 256'h3ef93ef941f8c2f96bf9f4f905fb92f8c9fed60ac20d510cf00b050ce00d1a0f;
// music[8253] = 256'he80e790fff0f4210b911c6126f1240128a11f1102611791049106810410f150f;
// music[8254] = 256'h370f610ed40e440f410f3211f612b9128f120813cf12e2124f15ef16cf156115;
// music[8255] = 256'h0015e3139b13511374137d131713b813ea135a149915e5159816441717173317;
// music[8256] = 256'h7617671838199019371afd19261ad3196317d516e0172e1874185318ec188a19;
// music[8257] = 256'h85198b1abb1a3c1a83198b1890195d19e417fa160d15af1591158914de155e0b;
// music[8258] = 256'h7100820cd9188d17bf1715184417a21874184e18fe180a19c719b61a031b811a;
// music[8259] = 256'h221a4f1af319071a171a8319d719391ab81abb1ba31b8a1b161c2c1c6d1cc91c;
// music[8260] = 256'hf71c321d571d9c1d511d1a1d851d011d001d1d1e801edb1e931ec01db11d781d;
// music[8261] = 256'h151eec1d691d4a1f9018bd092c05fe0684059e05a00582040c058704ff034804;
// music[8262] = 256'hcb03f60388040605d804a0036d0368035003dd0397038803de03470486058e05;
// music[8263] = 256'h1a051105f4032c0315033003b103050451041504fc03780458049004ee04ec04;
// music[8264] = 256'h16057f041a042a04f0032204f8034004cb0489045005c506a7090109c9fe4dfa;
// music[8265] = 256'he400ac0323065a0b800cf30def0efc0cfd0b180ac90769061004f401330088fe;
// music[8266] = 256'h9ffd95fe3a01d70179010202ef01df022b04cd04f80562061b068e06cd0adc10;
// music[8267] = 256'hbc10570f26120013d2122f146815611721198b1adc1b361d1f215424cf244926;
// music[8268] = 256'hcd27b228c8291c2a1f2b5d2cc72c912dbb2d6e2d8c2d062d4f2c892bd22be62d;
// music[8269] = 256'hc52ddf2b0e2b7b286a252f244e225621b2210321e2201421c220f320c7207620;
// music[8270] = 256'h5620f71f651f771eaa1d771bda188618c417ca169e155c138912840eb50e131d;
// music[8271] = 256'hdd2409206c1fd91ebe1bf81a6219ef181919f6171e18e5178c1775179f16aa16;
// music[8272] = 256'h0b16fd149d14be137213bd12a21151112b101d0f020eb40c550cdc0a62091009;
// music[8273] = 256'h62088f07b5052604f8034a0384024d017800380019ff4dffc1fe74fde5fd05fc;
// music[8274] = 256'h4dfc95fc60f36aefd9f43df404f34df56ff467f3f3f201f2eef1eaf0b9ef3cef;
// music[8275] = 256'h43ee5eedb3ec5bec3decc8eb48ebfdea4aebb8eb84eb76eb7feb16ebd3eab4ea;
// music[8276] = 256'h60ea0deaece9f0e9ebe9b4e995e9d4e90feaf2e9b9e9abe99de96be95ee928e9;
// music[8277] = 256'hcce8f9e8fde8b9e8d4e8e2e82be952e920e98de9b1e976e9c1e9f5e945eaacea;
// music[8278] = 256'he8ea32eb19eb37eba9eb49ec95ecadebf2eb35ec5bea10eb93ed26ee5eee56ee;
// music[8279] = 256'h34ef07f132f1c0f058f06ef032f076effcf0a5ec28e1a6dd1bdf22dd0cde8ce0;
// music[8280] = 256'hf4e044e10de154e1bde17ae1e2e1c1e1b1e1eae148e168e25be41ae478e389e3;
// music[8281] = 256'h96e3b1e3b9e3abe3bae3e2e3d5e309e47ee427e423e4a7e491e4fae481e4bde2;
// music[8282] = 256'hdbe28ee3b8e325e43ce31ae3b9e4e5e4a5e408e51de53ae518e565e542e6b1e6;
// music[8283] = 256'h1de7cee6a1e55de51de662e61ce62de60ee531e4e1e472e3ede732f662fc12f9;
// music[8284] = 256'h51f938fab7f921fa2efadffa10fbd5faa9fbe5fb38fc44fc74fb79fb67fb93fb;
// music[8285] = 256'h40fc48fc96fcb7fca6fcecfcfdfca1fd4afecefe6aff26ff2cff2effe2fe4eff;
// music[8286] = 256'h1bff26ff85fff3fe28ff86fffeffc1005a008f0092007000ac01f500f7017e02;
// music[8287] = 256'h46f7b6eb9beb77ec9beb86eca8ec2dedd5ed27ed4eed65ed32ec75eb9aebcfeb;
// music[8288] = 256'habebd3eb7fecd4ec3ced30eee9ee21ef79ef1cf052f03af04df057f066f087f0;
// music[8289] = 256'hbaf0c0f0b0f017f14ff16af182f1cdf07ff01ff1a0f108f23af259f2a6f280f2;
// music[8290] = 256'h6ef213f398f3d8f303f4def3f4f33ef444f46ff4e7f48cf5fdf5daf5bdf5d0f5;
// music[8291] = 256'hc9f50af66cf65af673f6a3f693f6eaf786f978f997f9c8f9cdf994fa3efa6ffa;
// music[8292] = 256'h93fc0afd59fc00fc3cfbe3faabfa7afa4afab3f938fac7fbadfc78fc48fc7ffc;
// music[8293] = 256'h87fcf6fc19fdd1fc67fcadfba5fb7efbfafbf3fc24fd42ff47001fff2aff94fe;
// music[8294] = 256'hb8fe12ff54fe99fef6fda0fdd8fd5bfd41fe30fea6fdb8fe8bffbeff65ffabff;
// music[8295] = 256'h2700d4ff180049ff61fdabfdeefebdfefdfe9cff5200ed00ebff88053510f112;
// music[8296] = 256'h02138f13de122114ba133e13be11b6109213921171169124be2625254a265f24;
// music[8297] = 256'h8a24a9242224b325cc262326ec249325f5252e261e2694247d253b251d244925;
// music[8298] = 256'hdb23ea230e26df25182689255925282795272b27b42749284d27ad2680270028;
// music[8299] = 256'h13286c26af25a12643263228ae2a0b2b9e2bf52a5b2a7b2ae62a132b21296f28;
// music[8300] = 256'hf427a327cd287d27ca265e278727c427ef269b2709274b264926d3232a26d123;
// music[8301] = 256'hb1133208ad099d097cfe6cf6eaf6e3f5b1f62ef7fdf51cf7e9f619f839f962f8;
// music[8302] = 256'h8bf9e6f8edf7c2f8dff79cf7abf80ef8c6f765f7a7f65df81bf929f930fa53f9;
// music[8303] = 256'heef9ccf95af702f7cbf6f5f669f8baf814f95efaeafa53fae4f83ff774fad9fe;
// music[8304] = 256'h76fe71fd7dfdf50095049c01f6fe6301e90552077d047d0117fe81f967f606f6;
// music[8305] = 256'h57f583f791fd3dfc53f2d3e606e55bee47f1cce8addc5ade4af3dd02d7037201;
// music[8306] = 256'hba08f415271136fc5df01cf5b4f953f268e075cdd4d367f23a099f11e311600d;
// music[8307] = 256'h1a0ae1098a09d607e6075108f6041f04c10da116ca11d70811094615a320621c;
// music[8308] = 256'ha00c4802c50a4019a819850ab7f1fde0bde30cf72e15952cf72e8d1dd906acfa;
// music[8309] = 256'hc2fd761194256b24b10f40f713ec63eceeee64f77cffb001b5051c0ebe17c618;
// music[8310] = 256'h9b0ef207f20c53141912d50729003f08a019c41d1021932819215e1a481b9f18;
// music[8311] = 256'hff17371dc227773105341a2c791eda1c7c26e12cd3303b401155176326686a5b;
// music[8312] = 256'hec4e8e50ef58bf6e9b7bff72505ef146ea420a406d319e20f70557f637fa35fa;
// music[8313] = 256'h65f362fa2f104c1ada15da0549ef79e62be8e9eaacee8ff5b6f75ded0eebc3f6;
// music[8314] = 256'h3a01dc092814e61cca20f921e824392cb4362d4356462a3db33fda40262b2516;
// music[8315] = 256'h3012c3187318c714271b6c1c191c9e252c2e9c2c9e240422c425da2a852ad220;
// music[8316] = 256'h111db123922965308e387736642bac1dd510fe08b105310c9b120b101d121918;
// music[8317] = 256'hed2ad244764f6751ad48213a7e283a09fbee9be126db8ad266c6b3cad3e4bb09;
// music[8318] = 256'h9e1d6819f61b9625cf25011dda17fa206f2ee531712db62fe539e4443f4e7151;
// music[8319] = 256'h5752ab50bf4bb6478245e64c7c5958612b632a612161665fb45f8d6636695c5e;
// music[8320] = 256'h4a476342ec554b5ebe5c945f36637f636b59bf4d384a945420683469b7611866;
// music[8321] = 256'h9b66b060855cc15fbc69406e3968d5574f4ae6448b3d993287216917d71ad219;
// music[8322] = 256'hff1925249f2acd241418df0a1b082f19eb29f222110e130ad21b5f272d277325;
// music[8323] = 256'h03227a15430e33241b2b450c36f95604471bac1fd813110e10092d0d5017e320;
// music[8324] = 256'h152b4b2bac2a0d23c60e2102e5fdc8036d0f3713b913a6134f0c75081814a924;
// music[8325] = 256'h1e335232bb1ae90d36181520291b8f1b862ba53c3d470e4ffc51ec40c61f920b;
// music[8326] = 256'hff06680ae1188a36d04cad440d415b4bc3471f362522b021bf2b65301039ac39;
// music[8327] = 256'h5831ee294b22c11e4521162cb03b8544c942fa40433cbe26cf13771512243833;
// music[8328] = 256'hac31631a7406520f5f28c63ad8389021e711cc167026a833322ee817e205650e;
// music[8329] = 256'h3b22bd27b226fc22a120c420fd1ab913570f4908ce003e0671108312e011ba0b;
// music[8330] = 256'hcf08610e6b11f60703eef8d79ed427e0e5ecadea80e682e7e0e997ee96ee97ea;
// music[8331] = 256'hdceb3df573fae2f67eef51e3cfe366f0cdf5b0f1c3e537e7c8fb3407ce05c105;
// music[8332] = 256'h030f871f4a29e221900ccdfd0704910dcb0785fb45fdd40f12176e0393f057f8;
// music[8333] = 256'h960d54159c11ba0fd9113517521169ff5ff657f60cfa6100200171febcfc12f7;
// music[8334] = 256'hcff152f115f6e1ff2efb39e5e5d965e45df2d3eca2e5f4ec11f568fdb3f9e1ed;
// music[8335] = 256'h86f0b2faaf00c7f592e94de9c0e59eee52fae4f441f1a7f6fb05ba1053101516;
// music[8336] = 256'h351a5a1b7f1ba914aa14331a081e50223122082600292f219e1c3316500810fc;
// music[8337] = 256'h2ef4d3f075ecc8fbda1bf423141e4f17040ec60be20f301c131f13188310a2f9;
// music[8338] = 256'h79eccff634082816040a9ff42ae712de51eb66f895efe5e8a2e86cef92fb4bfe;
// music[8339] = 256'h97f95ef153e9b6e2fbdc1ae016dc04cbd5c58ecd03d2b4ca6dbf35bc2ec5f9dd;
// music[8340] = 256'h7fee02e7b5df30e40bed36f285f0b1e5f4d1e2c544c5eac67bca33cb97c63bc3;
// music[8341] = 256'h5cc77ccf73ce3ad33eeb5bf63ef1dcf020eec4ed20ef2bee3bee01ec61efe5e3;
// music[8342] = 256'hadc938c63bc75bc424c8edc779c884c9abca3bc87cc407d490e8f2efedf062f0;
// music[8343] = 256'h8eeb57d88bc1a0c18dd751e825ebafec1fece7e734e6b0e65fe3d2d4b6c5dbc7;
// music[8344] = 256'hd0d34ede3fef7002050391f25ee799e5cadc4ecd77c7bfcfc1d967db6ce2a5ee;
// music[8345] = 256'h13efd8e84fe70cec63e497cf03ceb7e144f5a9f3ece1dfdaf1de33e0e3d290c9;
// music[8346] = 256'hbadd8ef5ccfce7fd1dfd14ecd7cdc5c496d485de33d99cdecef67c0439034a01;
// music[8347] = 256'h6cffddee73d5a0cf90d84ce7dcfa390e6f2275262d217722ed190d059bf817fc;
// music[8348] = 256'he0fb01f766ffd609540823041c0e0a1cae1d68144505c307631fdc2e07255a08;
// music[8349] = 256'h79f788ff9914f622c8172400a5f48000ee1a4628c51b2c0330f77104051c1121;
// music[8350] = 256'h660e66f5a2ec4bfe260740f71fe439cefbc4a0d58ceb67f2b6eb58edade9bfce;
// music[8351] = 256'h98bb5eb929b604b7d9bc31bcf2b7a7b33ab1fbb420b7c6b514b2c1aec2b132b4;
// music[8352] = 256'h92b5d1b724b80bb8b8b6e8b7f7b97cbb8ebdb5bbefb997ba42bbdfbb54bb74bb;
// music[8353] = 256'haebb50bc4ebfadbf20bf79cf1ae6a5e4b5d02fbd1abdb5d304e2aae157e13fe2;
// music[8354] = 256'h48e114df0add0cd83fd73edc30dc4bdb6adcfbdbced955d7a0d290cc9cca3fca;
// music[8355] = 256'h86cb2bcd3bcd6dcf61cd32c9c7c884cb2bcb70c6b4c907cb19cc5ad11abec1a7;
//     end
endmodule