module cos (input  logic        Clk,
            input  logic  [9:0] angle,
            output logic [20:0] answer);
    
    reg signed [10:0] cosine [0:1023];
    logic signed [10:0] answer_10;

    assign answer = {{10{answer_10[10]}}, answer_10};
    always_ff @ (posedge Clk) begin
        answer_10 <= cosine[angle];
    end

    initial begin
        cosine[0] = 11'sd1023;
        cosine[1] = 11'sd1022;
        cosine[2] = 11'sd1022;
        cosine[3] = 11'sd1022;
        cosine[4] = 11'sd1022;
        cosine[5] = 11'sd1022;
        cosine[6] = 11'sd1022;
        cosine[7] = 11'sd1022;
        cosine[8] = 11'sd1021;
        cosine[9] = 11'sd1021;
        cosine[10] = 11'sd1021;
        cosine[11] = 11'sd1020;
        cosine[12] = 11'sd1020;
        cosine[13] = 11'sd1019;
        cosine[14] = 11'sd1019;
        cosine[15] = 11'sd1018;
        cosine[16] = 11'sd1018;
        cosine[17] = 11'sd1017;
        cosine[18] = 11'sd1016;
        cosine[19] = 11'sd1016;
        cosine[20] = 11'sd1015;
        cosine[21] = 11'sd1014;
        cosine[22] = 11'sd1013;
        cosine[23] = 11'sd1012;
        cosine[24] = 11'sd1011;
        cosine[25] = 11'sd1010;
        cosine[26] = 11'sd1010;
        cosine[27] = 11'sd1008;
        cosine[28] = 11'sd1007;
        cosine[29] = 11'sd1006;
        cosine[30] = 11'sd1005;
        cosine[31] = 11'sd1004;
        cosine[32] = 11'sd1003;
        cosine[33] = 11'sd1002;
        cosine[34] = 11'sd1000;
        cosine[35] = 11'sd999;
        cosine[36] = 11'sd998;
        cosine[37] = 11'sd996;
        cosine[38] = 11'sd995;
        cosine[39] = 11'sd993;
        cosine[40] = 11'sd992;
        cosine[41] = 11'sd990;
        cosine[42] = 11'sd989;
        cosine[43] = 11'sd987;
        cosine[44] = 11'sd985;
        cosine[45] = 11'sd984;
        cosine[46] = 11'sd982;
        cosine[47] = 11'sd980;
        cosine[48] = 11'sd978;
        cosine[49] = 11'sd977;
        cosine[50] = 11'sd975;
        cosine[51] = 11'sd973;
        cosine[52] = 11'sd971;
        cosine[53] = 11'sd969;
        cosine[54] = 11'sd967;
        cosine[55] = 11'sd965;
        cosine[56] = 11'sd963;
        cosine[57] = 11'sd961;
        cosine[58] = 11'sd958;
        cosine[59] = 11'sd956;
        cosine[60] = 11'sd954;
        cosine[61] = 11'sd952;
        cosine[62] = 11'sd949;
        cosine[63] = 11'sd947;
        cosine[64] = 11'sd945;
        cosine[65] = 11'sd942;
        cosine[66] = 11'sd940;
        cosine[67] = 11'sd937;
        cosine[68] = 11'sd935;
        cosine[69] = 11'sd932;
        cosine[70] = 11'sd930;
        cosine[71] = 11'sd927;
        cosine[72] = 11'sd924;
        cosine[73] = 11'sd922;
        cosine[74] = 11'sd919;
        cosine[75] = 11'sd916;
        cosine[76] = 11'sd913;
        cosine[77] = 11'sd910;
        cosine[78] = 11'sd908;
        cosine[79] = 11'sd905;
        cosine[80] = 11'sd902;
        cosine[81] = 11'sd899;
        cosine[82] = 11'sd896;
        cosine[83] = 11'sd893;
        cosine[84] = 11'sd890;
        cosine[85] = 11'sd886;
        cosine[86] = 11'sd883;
        cosine[87] = 11'sd880;
        cosine[88] = 11'sd877;
        cosine[89] = 11'sd874;
        cosine[90] = 11'sd870;
        cosine[91] = 11'sd867;
        cosine[92] = 11'sd864;
        cosine[93] = 11'sd860;
        cosine[94] = 11'sd857;
        cosine[95] = 11'sd854;
        cosine[96] = 11'sd850;
        cosine[97] = 11'sd847;
        cosine[98] = 11'sd843;
        cosine[99] = 11'sd839;
        cosine[100] = 11'sd836;
        cosine[101] = 11'sd832;
        cosine[102] = 11'sd829;
        cosine[103] = 11'sd825;
        cosine[104] = 11'sd821;
        cosine[105] = 11'sd817;
        cosine[106] = 11'sd814;
        cosine[107] = 11'sd810;
        cosine[108] = 11'sd806;
        cosine[109] = 11'sd802;
        cosine[110] = 11'sd798;
        cosine[111] = 11'sd794;
        cosine[112] = 11'sd790;
        cosine[113] = 11'sd786;
        cosine[114] = 11'sd782;
        cosine[115] = 11'sd778;
        cosine[116] = 11'sd774;
        cosine[117] = 11'sd770;
        cosine[118] = 11'sd766;
        cosine[119] = 11'sd762;
        cosine[120] = 11'sd757;
        cosine[121] = 11'sd753;
        cosine[122] = 11'sd749;
        cosine[123] = 11'sd745;
        cosine[124] = 11'sd740;
        cosine[125] = 11'sd736;
        cosine[126] = 11'sd732;
        cosine[127] = 11'sd727;
        cosine[128] = 11'sd723;
        cosine[129] = 11'sd718;
        cosine[130] = 11'sd714;
        cosine[131] = 11'sd709;
        cosine[132] = 11'sd705;
        cosine[133] = 11'sd700;
        cosine[134] = 11'sd696;
        cosine[135] = 11'sd691;
        cosine[136] = 11'sd687;
        cosine[137] = 11'sd682;
        cosine[138] = 11'sd677;
        cosine[139] = 11'sd672;
        cosine[140] = 11'sd668;
        cosine[141] = 11'sd663;
        cosine[142] = 11'sd658;
        cosine[143] = 11'sd653;
        cosine[144] = 11'sd648;
        cosine[145] = 11'sd644;
        cosine[146] = 11'sd639;
        cosine[147] = 11'sd634;
        cosine[148] = 11'sd629;
        cosine[149] = 11'sd624;
        cosine[150] = 11'sd619;
        cosine[151] = 11'sd614;
        cosine[152] = 11'sd609;
        cosine[153] = 11'sd604;
        cosine[154] = 11'sd599;
        cosine[155] = 11'sd594;
        cosine[156] = 11'sd589;
        cosine[157] = 11'sd583;
        cosine[158] = 11'sd578;
        cosine[159] = 11'sd573;
        cosine[160] = 11'sd568;
        cosine[161] = 11'sd563;
        cosine[162] = 11'sd557;
        cosine[163] = 11'sd552;
        cosine[164] = 11'sd547;
        cosine[165] = 11'sd541;
        cosine[166] = 11'sd536;
        cosine[167] = 11'sd531;
        cosine[168] = 11'sd525;
        cosine[169] = 11'sd520;
        cosine[170] = 11'sd515;
        cosine[171] = 11'sd509;
        cosine[172] = 11'sd504;
        cosine[173] = 11'sd498;
        cosine[174] = 11'sd493;
        cosine[175] = 11'sd487;
        cosine[176] = 11'sd482;
        cosine[177] = 11'sd476;
        cosine[178] = 11'sd471;
        cosine[179] = 11'sd465;
        cosine[180] = 11'sd459;
        cosine[181] = 11'sd454;
        cosine[182] = 11'sd448;
        cosine[183] = 11'sd443;
        cosine[184] = 11'sd437;
        cosine[185] = 11'sd431;
        cosine[186] = 11'sd426;
        cosine[187] = 11'sd420;
        cosine[188] = 11'sd414;
        cosine[189] = 11'sd408;
        cosine[190] = 11'sd403;
        cosine[191] = 11'sd397;
        cosine[192] = 11'sd391;
        cosine[193] = 11'sd385;
        cosine[194] = 11'sd379;
        cosine[195] = 11'sd374;
        cosine[196] = 11'sd368;
        cosine[197] = 11'sd362;
        cosine[198] = 11'sd356;
        cosine[199] = 11'sd350;
        cosine[200] = 11'sd344;
        cosine[201] = 11'sd338;
        cosine[202] = 11'sd332;
        cosine[203] = 11'sd326;
        cosine[204] = 11'sd320;
        cosine[205] = 11'sd314;
        cosine[206] = 11'sd308;
        cosine[207] = 11'sd302;
        cosine[208] = 11'sd296;
        cosine[209] = 11'sd290;
        cosine[210] = 11'sd284;
        cosine[211] = 11'sd278;
        cosine[212] = 11'sd272;
        cosine[213] = 11'sd266;
        cosine[214] = 11'sd260;
        cosine[215] = 11'sd254;
        cosine[216] = 11'sd248;
        cosine[217] = 11'sd242;
        cosine[218] = 11'sd236;
        cosine[219] = 11'sd230;
        cosine[220] = 11'sd224;
        cosine[221] = 11'sd218;
        cosine[222] = 11'sd211;
        cosine[223] = 11'sd205;
        cosine[224] = 11'sd199;
        cosine[225] = 11'sd193;
        cosine[226] = 11'sd187;
        cosine[227] = 11'sd181;
        cosine[228] = 11'sd174;
        cosine[229] = 11'sd168;
        cosine[230] = 11'sd162;
        cosine[231] = 11'sd156;
        cosine[232] = 11'sd150;
        cosine[233] = 11'sd143;
        cosine[234] = 11'sd137;
        cosine[235] = 11'sd131;
        cosine[236] = 11'sd125;
        cosine[237] = 11'sd118;
        cosine[238] = 11'sd112;
        cosine[239] = 11'sd106;
        cosine[240] = 11'sd100;
        cosine[241] = 11'sd94;
        cosine[242] = 11'sd87;
        cosine[243] = 11'sd81;
        cosine[244] = 11'sd75;
        cosine[245] = 11'sd68;
        cosine[246] = 11'sd62;
        cosine[247] = 11'sd56;
        cosine[248] = 11'sd50;
        cosine[249] = 11'sd43;
        cosine[250] = 11'sd37;
        cosine[251] = 11'sd31;
        cosine[252] = 11'sd25;
        cosine[253] = 11'sd18;
        cosine[254] = 11'sd12;
        cosine[255] = 11'sd6;
        cosine[256] = 11'sd0;
        cosine[257] = -11'sd6;
        cosine[258] = -11'sd12;
        cosine[259] = -11'sd18;
        cosine[260] = -11'sd25;
        cosine[261] = -11'sd31;
        cosine[262] = -11'sd37;
        cosine[263] = -11'sd43;
        cosine[264] = -11'sd50;
        cosine[265] = -11'sd56;
        cosine[266] = -11'sd62;
        cosine[267] = -11'sd68;
        cosine[268] = -11'sd75;
        cosine[269] = -11'sd81;
        cosine[270] = -11'sd87;
        cosine[271] = -11'sd94;
        cosine[272] = -11'sd100;
        cosine[273] = -11'sd106;
        cosine[274] = -11'sd112;
        cosine[275] = -11'sd118;
        cosine[276] = -11'sd125;
        cosine[277] = -11'sd131;
        cosine[278] = -11'sd137;
        cosine[279] = -11'sd143;
        cosine[280] = -11'sd150;
        cosine[281] = -11'sd156;
        cosine[282] = -11'sd162;
        cosine[283] = -11'sd168;
        cosine[284] = -11'sd174;
        cosine[285] = -11'sd181;
        cosine[286] = -11'sd187;
        cosine[287] = -11'sd193;
        cosine[288] = -11'sd199;
        cosine[289] = -11'sd205;
        cosine[290] = -11'sd211;
        cosine[291] = -11'sd218;
        cosine[292] = -11'sd224;
        cosine[293] = -11'sd230;
        cosine[294] = -11'sd236;
        cosine[295] = -11'sd242;
        cosine[296] = -11'sd248;
        cosine[297] = -11'sd254;
        cosine[298] = -11'sd260;
        cosine[299] = -11'sd266;
        cosine[300] = -11'sd272;
        cosine[301] = -11'sd278;
        cosine[302] = -11'sd284;
        cosine[303] = -11'sd290;
        cosine[304] = -11'sd296;
        cosine[305] = -11'sd302;
        cosine[306] = -11'sd308;
        cosine[307] = -11'sd314;
        cosine[308] = -11'sd320;
        cosine[309] = -11'sd326;
        cosine[310] = -11'sd332;
        cosine[311] = -11'sd338;
        cosine[312] = -11'sd344;
        cosine[313] = -11'sd350;
        cosine[314] = -11'sd356;
        cosine[315] = -11'sd362;
        cosine[316] = -11'sd368;
        cosine[317] = -11'sd374;
        cosine[318] = -11'sd379;
        cosine[319] = -11'sd385;
        cosine[320] = -11'sd391;
        cosine[321] = -11'sd397;
        cosine[322] = -11'sd403;
        cosine[323] = -11'sd408;
        cosine[324] = -11'sd414;
        cosine[325] = -11'sd420;
        cosine[326] = -11'sd426;
        cosine[327] = -11'sd431;
        cosine[328] = -11'sd437;
        cosine[329] = -11'sd443;
        cosine[330] = -11'sd448;
        cosine[331] = -11'sd454;
        cosine[332] = -11'sd459;
        cosine[333] = -11'sd465;
        cosine[334] = -11'sd471;
        cosine[335] = -11'sd476;
        cosine[336] = -11'sd482;
        cosine[337] = -11'sd487;
        cosine[338] = -11'sd493;
        cosine[339] = -11'sd498;
        cosine[340] = -11'sd504;
        cosine[341] = -11'sd509;
        cosine[342] = -11'sd515;
        cosine[343] = -11'sd520;
        cosine[344] = -11'sd525;
        cosine[345] = -11'sd531;
        cosine[346] = -11'sd536;
        cosine[347] = -11'sd541;
        cosine[348] = -11'sd547;
        cosine[349] = -11'sd552;
        cosine[350] = -11'sd557;
        cosine[351] = -11'sd563;
        cosine[352] = -11'sd568;
        cosine[353] = -11'sd573;
        cosine[354] = -11'sd578;
        cosine[355] = -11'sd583;
        cosine[356] = -11'sd589;
        cosine[357] = -11'sd594;
        cosine[358] = -11'sd599;
        cosine[359] = -11'sd604;
        cosine[360] = -11'sd609;
        cosine[361] = -11'sd614;
        cosine[362] = -11'sd619;
        cosine[363] = -11'sd624;
        cosine[364] = -11'sd629;
        cosine[365] = -11'sd634;
        cosine[366] = -11'sd639;
        cosine[367] = -11'sd644;
        cosine[368] = -11'sd648;
        cosine[369] = -11'sd653;
        cosine[370] = -11'sd658;
        cosine[371] = -11'sd663;
        cosine[372] = -11'sd668;
        cosine[373] = -11'sd672;
        cosine[374] = -11'sd677;
        cosine[375] = -11'sd682;
        cosine[376] = -11'sd687;
        cosine[377] = -11'sd691;
        cosine[378] = -11'sd696;
        cosine[379] = -11'sd700;
        cosine[380] = -11'sd705;
        cosine[381] = -11'sd709;
        cosine[382] = -11'sd714;
        cosine[383] = -11'sd718;
        cosine[384] = -11'sd723;
        cosine[385] = -11'sd727;
        cosine[386] = -11'sd732;
        cosine[387] = -11'sd736;
        cosine[388] = -11'sd740;
        cosine[389] = -11'sd745;
        cosine[390] = -11'sd749;
        cosine[391] = -11'sd753;
        cosine[392] = -11'sd757;
        cosine[393] = -11'sd762;
        cosine[394] = -11'sd766;
        cosine[395] = -11'sd770;
        cosine[396] = -11'sd774;
        cosine[397] = -11'sd778;
        cosine[398] = -11'sd782;
        cosine[399] = -11'sd786;
        cosine[400] = -11'sd790;
        cosine[401] = -11'sd794;
        cosine[402] = -11'sd798;
        cosine[403] = -11'sd802;
        cosine[404] = -11'sd806;
        cosine[405] = -11'sd810;
        cosine[406] = -11'sd814;
        cosine[407] = -11'sd817;
        cosine[408] = -11'sd821;
        cosine[409] = -11'sd825;
        cosine[410] = -11'sd829;
        cosine[411] = -11'sd832;
        cosine[412] = -11'sd836;
        cosine[413] = -11'sd839;
        cosine[414] = -11'sd843;
        cosine[415] = -11'sd847;
        cosine[416] = -11'sd850;
        cosine[417] = -11'sd854;
        cosine[418] = -11'sd857;
        cosine[419] = -11'sd860;
        cosine[420] = -11'sd864;
        cosine[421] = -11'sd867;
        cosine[422] = -11'sd870;
        cosine[423] = -11'sd874;
        cosine[424] = -11'sd877;
        cosine[425] = -11'sd880;
        cosine[426] = -11'sd883;
        cosine[427] = -11'sd886;
        cosine[428] = -11'sd890;
        cosine[429] = -11'sd893;
        cosine[430] = -11'sd896;
        cosine[431] = -11'sd899;
        cosine[432] = -11'sd902;
        cosine[433] = -11'sd905;
        cosine[434] = -11'sd908;
        cosine[435] = -11'sd910;
        cosine[436] = -11'sd913;
        cosine[437] = -11'sd916;
        cosine[438] = -11'sd919;
        cosine[439] = -11'sd922;
        cosine[440] = -11'sd924;
        cosine[441] = -11'sd927;
        cosine[442] = -11'sd930;
        cosine[443] = -11'sd932;
        cosine[444] = -11'sd935;
        cosine[445] = -11'sd937;
        cosine[446] = -11'sd940;
        cosine[447] = -11'sd942;
        cosine[448] = -11'sd945;
        cosine[449] = -11'sd947;
        cosine[450] = -11'sd949;
        cosine[451] = -11'sd952;
        cosine[452] = -11'sd954;
        cosine[453] = -11'sd956;
        cosine[454] = -11'sd958;
        cosine[455] = -11'sd961;
        cosine[456] = -11'sd963;
        cosine[457] = -11'sd965;
        cosine[458] = -11'sd967;
        cosine[459] = -11'sd969;
        cosine[460] = -11'sd971;
        cosine[461] = -11'sd973;
        cosine[462] = -11'sd975;
        cosine[463] = -11'sd977;
        cosine[464] = -11'sd978;
        cosine[465] = -11'sd980;
        cosine[466] = -11'sd982;
        cosine[467] = -11'sd984;
        cosine[468] = -11'sd985;
        cosine[469] = -11'sd987;
        cosine[470] = -11'sd989;
        cosine[471] = -11'sd990;
        cosine[472] = -11'sd992;
        cosine[473] = -11'sd993;
        cosine[474] = -11'sd995;
        cosine[475] = -11'sd996;
        cosine[476] = -11'sd998;
        cosine[477] = -11'sd999;
        cosine[478] = -11'sd1000;
        cosine[479] = -11'sd1002;
        cosine[480] = -11'sd1003;
        cosine[481] = -11'sd1004;
        cosine[482] = -11'sd1005;
        cosine[483] = -11'sd1006;
        cosine[484] = -11'sd1007;
        cosine[485] = -11'sd1008;
        cosine[486] = -11'sd1010;
        cosine[487] = -11'sd1010;
        cosine[488] = -11'sd1011;
        cosine[489] = -11'sd1012;
        cosine[490] = -11'sd1013;
        cosine[491] = -11'sd1014;
        cosine[492] = -11'sd1015;
        cosine[493] = -11'sd1016;
        cosine[494] = -11'sd1016;
        cosine[495] = -11'sd1017;
        cosine[496] = -11'sd1018;
        cosine[497] = -11'sd1018;
        cosine[498] = -11'sd1019;
        cosine[499] = -11'sd1019;
        cosine[500] = -11'sd1020;
        cosine[501] = -11'sd1020;
        cosine[502] = -11'sd1021;
        cosine[503] = -11'sd1021;
        cosine[504] = -11'sd1021;
        cosine[505] = -11'sd1022;
        cosine[506] = -11'sd1022;
        cosine[507] = -11'sd1022;
        cosine[508] = -11'sd1022;
        cosine[509] = -11'sd1022;
        cosine[510] = -11'sd1022;
        cosine[511] = -11'sd1022;
        cosine[512] = -11'sd1023;
        cosine[513] = -11'sd1022;
        cosine[514] = -11'sd1022;
        cosine[515] = -11'sd1022;
        cosine[516] = -11'sd1022;
        cosine[517] = -11'sd1022;
        cosine[518] = -11'sd1022;
        cosine[519] = -11'sd1022;
        cosine[520] = -11'sd1021;
        cosine[521] = -11'sd1021;
        cosine[522] = -11'sd1021;
        cosine[523] = -11'sd1020;
        cosine[524] = -11'sd1020;
        cosine[525] = -11'sd1019;
        cosine[526] = -11'sd1019;
        cosine[527] = -11'sd1018;
        cosine[528] = -11'sd1018;
        cosine[529] = -11'sd1017;
        cosine[530] = -11'sd1016;
        cosine[531] = -11'sd1016;
        cosine[532] = -11'sd1015;
        cosine[533] = -11'sd1014;
        cosine[534] = -11'sd1013;
        cosine[535] = -11'sd1012;
        cosine[536] = -11'sd1011;
        cosine[537] = -11'sd1010;
        cosine[538] = -11'sd1010;
        cosine[539] = -11'sd1008;
        cosine[540] = -11'sd1007;
        cosine[541] = -11'sd1006;
        cosine[542] = -11'sd1005;
        cosine[543] = -11'sd1004;
        cosine[544] = -11'sd1003;
        cosine[545] = -11'sd1002;
        cosine[546] = -11'sd1000;
        cosine[547] = -11'sd999;
        cosine[548] = -11'sd998;
        cosine[549] = -11'sd996;
        cosine[550] = -11'sd995;
        cosine[551] = -11'sd993;
        cosine[552] = -11'sd992;
        cosine[553] = -11'sd990;
        cosine[554] = -11'sd989;
        cosine[555] = -11'sd987;
        cosine[556] = -11'sd985;
        cosine[557] = -11'sd984;
        cosine[558] = -11'sd982;
        cosine[559] = -11'sd980;
        cosine[560] = -11'sd978;
        cosine[561] = -11'sd977;
        cosine[562] = -11'sd975;
        cosine[563] = -11'sd973;
        cosine[564] = -11'sd971;
        cosine[565] = -11'sd969;
        cosine[566] = -11'sd967;
        cosine[567] = -11'sd965;
        cosine[568] = -11'sd963;
        cosine[569] = -11'sd961;
        cosine[570] = -11'sd958;
        cosine[571] = -11'sd956;
        cosine[572] = -11'sd954;
        cosine[573] = -11'sd952;
        cosine[574] = -11'sd949;
        cosine[575] = -11'sd947;
        cosine[576] = -11'sd945;
        cosine[577] = -11'sd942;
        cosine[578] = -11'sd940;
        cosine[579] = -11'sd937;
        cosine[580] = -11'sd935;
        cosine[581] = -11'sd932;
        cosine[582] = -11'sd930;
        cosine[583] = -11'sd927;
        cosine[584] = -11'sd924;
        cosine[585] = -11'sd922;
        cosine[586] = -11'sd919;
        cosine[587] = -11'sd916;
        cosine[588] = -11'sd913;
        cosine[589] = -11'sd910;
        cosine[590] = -11'sd908;
        cosine[591] = -11'sd905;
        cosine[592] = -11'sd902;
        cosine[593] = -11'sd899;
        cosine[594] = -11'sd896;
        cosine[595] = -11'sd893;
        cosine[596] = -11'sd890;
        cosine[597] = -11'sd886;
        cosine[598] = -11'sd883;
        cosine[599] = -11'sd880;
        cosine[600] = -11'sd877;
        cosine[601] = -11'sd874;
        cosine[602] = -11'sd870;
        cosine[603] = -11'sd867;
        cosine[604] = -11'sd864;
        cosine[605] = -11'sd860;
        cosine[606] = -11'sd857;
        cosine[607] = -11'sd854;
        cosine[608] = -11'sd850;
        cosine[609] = -11'sd847;
        cosine[610] = -11'sd843;
        cosine[611] = -11'sd839;
        cosine[612] = -11'sd836;
        cosine[613] = -11'sd832;
        cosine[614] = -11'sd829;
        cosine[615] = -11'sd825;
        cosine[616] = -11'sd821;
        cosine[617] = -11'sd817;
        cosine[618] = -11'sd814;
        cosine[619] = -11'sd810;
        cosine[620] = -11'sd806;
        cosine[621] = -11'sd802;
        cosine[622] = -11'sd798;
        cosine[623] = -11'sd794;
        cosine[624] = -11'sd790;
        cosine[625] = -11'sd786;
        cosine[626] = -11'sd782;
        cosine[627] = -11'sd778;
        cosine[628] = -11'sd774;
        cosine[629] = -11'sd770;
        cosine[630] = -11'sd766;
        cosine[631] = -11'sd762;
        cosine[632] = -11'sd757;
        cosine[633] = -11'sd753;
        cosine[634] = -11'sd749;
        cosine[635] = -11'sd745;
        cosine[636] = -11'sd740;
        cosine[637] = -11'sd736;
        cosine[638] = -11'sd732;
        cosine[639] = -11'sd727;
        cosine[640] = -11'sd723;
        cosine[641] = -11'sd718;
        cosine[642] = -11'sd714;
        cosine[643] = -11'sd709;
        cosine[644] = -11'sd705;
        cosine[645] = -11'sd700;
        cosine[646] = -11'sd696;
        cosine[647] = -11'sd691;
        cosine[648] = -11'sd687;
        cosine[649] = -11'sd682;
        cosine[650] = -11'sd677;
        cosine[651] = -11'sd672;
        cosine[652] = -11'sd668;
        cosine[653] = -11'sd663;
        cosine[654] = -11'sd658;
        cosine[655] = -11'sd653;
        cosine[656] = -11'sd648;
        cosine[657] = -11'sd644;
        cosine[658] = -11'sd639;
        cosine[659] = -11'sd634;
        cosine[660] = -11'sd629;
        cosine[661] = -11'sd624;
        cosine[662] = -11'sd619;
        cosine[663] = -11'sd614;
        cosine[664] = -11'sd609;
        cosine[665] = -11'sd604;
        cosine[666] = -11'sd599;
        cosine[667] = -11'sd594;
        cosine[668] = -11'sd589;
        cosine[669] = -11'sd583;
        cosine[670] = -11'sd578;
        cosine[671] = -11'sd573;
        cosine[672] = -11'sd568;
        cosine[673] = -11'sd563;
        cosine[674] = -11'sd557;
        cosine[675] = -11'sd552;
        cosine[676] = -11'sd547;
        cosine[677] = -11'sd541;
        cosine[678] = -11'sd536;
        cosine[679] = -11'sd531;
        cosine[680] = -11'sd525;
        cosine[681] = -11'sd520;
        cosine[682] = -11'sd515;
        cosine[683] = -11'sd509;
        cosine[684] = -11'sd504;
        cosine[685] = -11'sd498;
        cosine[686] = -11'sd493;
        cosine[687] = -11'sd487;
        cosine[688] = -11'sd482;
        cosine[689] = -11'sd476;
        cosine[690] = -11'sd471;
        cosine[691] = -11'sd465;
        cosine[692] = -11'sd459;
        cosine[693] = -11'sd454;
        cosine[694] = -11'sd448;
        cosine[695] = -11'sd443;
        cosine[696] = -11'sd437;
        cosine[697] = -11'sd431;
        cosine[698] = -11'sd426;
        cosine[699] = -11'sd420;
        cosine[700] = -11'sd414;
        cosine[701] = -11'sd408;
        cosine[702] = -11'sd403;
        cosine[703] = -11'sd397;
        cosine[704] = -11'sd391;
        cosine[705] = -11'sd385;
        cosine[706] = -11'sd379;
        cosine[707] = -11'sd374;
        cosine[708] = -11'sd368;
        cosine[709] = -11'sd362;
        cosine[710] = -11'sd356;
        cosine[711] = -11'sd350;
        cosine[712] = -11'sd344;
        cosine[713] = -11'sd338;
        cosine[714] = -11'sd332;
        cosine[715] = -11'sd326;
        cosine[716] = -11'sd320;
        cosine[717] = -11'sd314;
        cosine[718] = -11'sd308;
        cosine[719] = -11'sd302;
        cosine[720] = -11'sd296;
        cosine[721] = -11'sd290;
        cosine[722] = -11'sd284;
        cosine[723] = -11'sd278;
        cosine[724] = -11'sd272;
        cosine[725] = -11'sd266;
        cosine[726] = -11'sd260;
        cosine[727] = -11'sd254;
        cosine[728] = -11'sd248;
        cosine[729] = -11'sd242;
        cosine[730] = -11'sd236;
        cosine[731] = -11'sd230;
        cosine[732] = -11'sd224;
        cosine[733] = -11'sd218;
        cosine[734] = -11'sd211;
        cosine[735] = -11'sd205;
        cosine[736] = -11'sd199;
        cosine[737] = -11'sd193;
        cosine[738] = -11'sd187;
        cosine[739] = -11'sd181;
        cosine[740] = -11'sd174;
        cosine[741] = -11'sd168;
        cosine[742] = -11'sd162;
        cosine[743] = -11'sd156;
        cosine[744] = -11'sd150;
        cosine[745] = -11'sd143;
        cosine[746] = -11'sd137;
        cosine[747] = -11'sd131;
        cosine[748] = -11'sd125;
        cosine[749] = -11'sd118;
        cosine[750] = -11'sd112;
        cosine[751] = -11'sd106;
        cosine[752] = -11'sd100;
        cosine[753] = -11'sd94;
        cosine[754] = -11'sd87;
        cosine[755] = -11'sd81;
        cosine[756] = -11'sd75;
        cosine[757] = -11'sd68;
        cosine[758] = -11'sd62;
        cosine[759] = -11'sd56;
        cosine[760] = -11'sd50;
        cosine[761] = -11'sd43;
        cosine[762] = -11'sd37;
        cosine[763] = -11'sd31;
        cosine[764] = -11'sd25;
        cosine[765] = -11'sd18;
        cosine[766] = -11'sd12;
        cosine[767] = -11'sd6;
        cosine[768] = 11'sd0;
        cosine[769] = 11'sd6;
        cosine[770] = 11'sd12;
        cosine[771] = 11'sd18;
        cosine[772] = 11'sd25;
        cosine[773] = 11'sd31;
        cosine[774] = 11'sd37;
        cosine[775] = 11'sd43;
        cosine[776] = 11'sd50;
        cosine[777] = 11'sd56;
        cosine[778] = 11'sd62;
        cosine[779] = 11'sd68;
        cosine[780] = 11'sd75;
        cosine[781] = 11'sd81;
        cosine[782] = 11'sd87;
        cosine[783] = 11'sd94;
        cosine[784] = 11'sd100;
        cosine[785] = 11'sd106;
        cosine[786] = 11'sd112;
        cosine[787] = 11'sd118;
        cosine[788] = 11'sd125;
        cosine[789] = 11'sd131;
        cosine[790] = 11'sd137;
        cosine[791] = 11'sd143;
        cosine[792] = 11'sd150;
        cosine[793] = 11'sd156;
        cosine[794] = 11'sd162;
        cosine[795] = 11'sd168;
        cosine[796] = 11'sd174;
        cosine[797] = 11'sd181;
        cosine[798] = 11'sd187;
        cosine[799] = 11'sd193;
        cosine[800] = 11'sd199;
        cosine[801] = 11'sd205;
        cosine[802] = 11'sd211;
        cosine[803] = 11'sd218;
        cosine[804] = 11'sd224;
        cosine[805] = 11'sd230;
        cosine[806] = 11'sd236;
        cosine[807] = 11'sd242;
        cosine[808] = 11'sd248;
        cosine[809] = 11'sd254;
        cosine[810] = 11'sd260;
        cosine[811] = 11'sd266;
        cosine[812] = 11'sd272;
        cosine[813] = 11'sd278;
        cosine[814] = 11'sd284;
        cosine[815] = 11'sd290;
        cosine[816] = 11'sd296;
        cosine[817] = 11'sd302;
        cosine[818] = 11'sd308;
        cosine[819] = 11'sd314;
        cosine[820] = 11'sd320;
        cosine[821] = 11'sd326;
        cosine[822] = 11'sd332;
        cosine[823] = 11'sd338;
        cosine[824] = 11'sd344;
        cosine[825] = 11'sd350;
        cosine[826] = 11'sd356;
        cosine[827] = 11'sd362;
        cosine[828] = 11'sd368;
        cosine[829] = 11'sd374;
        cosine[830] = 11'sd379;
        cosine[831] = 11'sd385;
        cosine[832] = 11'sd391;
        cosine[833] = 11'sd397;
        cosine[834] = 11'sd403;
        cosine[835] = 11'sd408;
        cosine[836] = 11'sd414;
        cosine[837] = 11'sd420;
        cosine[838] = 11'sd426;
        cosine[839] = 11'sd431;
        cosine[840] = 11'sd437;
        cosine[841] = 11'sd443;
        cosine[842] = 11'sd448;
        cosine[843] = 11'sd454;
        cosine[844] = 11'sd459;
        cosine[845] = 11'sd465;
        cosine[846] = 11'sd471;
        cosine[847] = 11'sd476;
        cosine[848] = 11'sd482;
        cosine[849] = 11'sd487;
        cosine[850] = 11'sd493;
        cosine[851] = 11'sd498;
        cosine[852] = 11'sd504;
        cosine[853] = 11'sd509;
        cosine[854] = 11'sd515;
        cosine[855] = 11'sd520;
        cosine[856] = 11'sd525;
        cosine[857] = 11'sd531;
        cosine[858] = 11'sd536;
        cosine[859] = 11'sd541;
        cosine[860] = 11'sd547;
        cosine[861] = 11'sd552;
        cosine[862] = 11'sd557;
        cosine[863] = 11'sd563;
        cosine[864] = 11'sd568;
        cosine[865] = 11'sd573;
        cosine[866] = 11'sd578;
        cosine[867] = 11'sd583;
        cosine[868] = 11'sd589;
        cosine[869] = 11'sd594;
        cosine[870] = 11'sd599;
        cosine[871] = 11'sd604;
        cosine[872] = 11'sd609;
        cosine[873] = 11'sd614;
        cosine[874] = 11'sd619;
        cosine[875] = 11'sd624;
        cosine[876] = 11'sd629;
        cosine[877] = 11'sd634;
        cosine[878] = 11'sd639;
        cosine[879] = 11'sd644;
        cosine[880] = 11'sd648;
        cosine[881] = 11'sd653;
        cosine[882] = 11'sd658;
        cosine[883] = 11'sd663;
        cosine[884] = 11'sd668;
        cosine[885] = 11'sd672;
        cosine[886] = 11'sd677;
        cosine[887] = 11'sd682;
        cosine[888] = 11'sd687;
        cosine[889] = 11'sd691;
        cosine[890] = 11'sd696;
        cosine[891] = 11'sd700;
        cosine[892] = 11'sd705;
        cosine[893] = 11'sd709;
        cosine[894] = 11'sd714;
        cosine[895] = 11'sd718;
        cosine[896] = 11'sd723;
        cosine[897] = 11'sd727;
        cosine[898] = 11'sd732;
        cosine[899] = 11'sd736;
        cosine[900] = 11'sd740;
        cosine[901] = 11'sd745;
        cosine[902] = 11'sd749;
        cosine[903] = 11'sd753;
        cosine[904] = 11'sd757;
        cosine[905] = 11'sd762;
        cosine[906] = 11'sd766;
        cosine[907] = 11'sd770;
        cosine[908] = 11'sd774;
        cosine[909] = 11'sd778;
        cosine[910] = 11'sd782;
        cosine[911] = 11'sd786;
        cosine[912] = 11'sd790;
        cosine[913] = 11'sd794;
        cosine[914] = 11'sd798;
        cosine[915] = 11'sd802;
        cosine[916] = 11'sd806;
        cosine[917] = 11'sd810;
        cosine[918] = 11'sd814;
        cosine[919] = 11'sd817;
        cosine[920] = 11'sd821;
        cosine[921] = 11'sd825;
        cosine[922] = 11'sd829;
        cosine[923] = 11'sd832;
        cosine[924] = 11'sd836;
        cosine[925] = 11'sd839;
        cosine[926] = 11'sd843;
        cosine[927] = 11'sd847;
        cosine[928] = 11'sd850;
        cosine[929] = 11'sd854;
        cosine[930] = 11'sd857;
        cosine[931] = 11'sd860;
        cosine[932] = 11'sd864;
        cosine[933] = 11'sd867;
        cosine[934] = 11'sd870;
        cosine[935] = 11'sd874;
        cosine[936] = 11'sd877;
        cosine[937] = 11'sd880;
        cosine[938] = 11'sd883;
        cosine[939] = 11'sd886;
        cosine[940] = 11'sd890;
        cosine[941] = 11'sd893;
        cosine[942] = 11'sd896;
        cosine[943] = 11'sd899;
        cosine[944] = 11'sd902;
        cosine[945] = 11'sd905;
        cosine[946] = 11'sd908;
        cosine[947] = 11'sd910;
        cosine[948] = 11'sd913;
        cosine[949] = 11'sd916;
        cosine[950] = 11'sd919;
        cosine[951] = 11'sd922;
        cosine[952] = 11'sd924;
        cosine[953] = 11'sd927;
        cosine[954] = 11'sd930;
        cosine[955] = 11'sd932;
        cosine[956] = 11'sd935;
        cosine[957] = 11'sd937;
        cosine[958] = 11'sd940;
        cosine[959] = 11'sd942;
        cosine[960] = 11'sd945;
        cosine[961] = 11'sd947;
        cosine[962] = 11'sd949;
        cosine[963] = 11'sd952;
        cosine[964] = 11'sd954;
        cosine[965] = 11'sd956;
        cosine[966] = 11'sd958;
        cosine[967] = 11'sd961;
        cosine[968] = 11'sd963;
        cosine[969] = 11'sd965;
        cosine[970] = 11'sd967;
        cosine[971] = 11'sd969;
        cosine[972] = 11'sd971;
        cosine[973] = 11'sd973;
        cosine[974] = 11'sd975;
        cosine[975] = 11'sd977;
        cosine[976] = 11'sd978;
        cosine[977] = 11'sd980;
        cosine[978] = 11'sd982;
        cosine[979] = 11'sd984;
        cosine[980] = 11'sd985;
        cosine[981] = 11'sd987;
        cosine[982] = 11'sd989;
        cosine[983] = 11'sd990;
        cosine[984] = 11'sd992;
        cosine[985] = 11'sd993;
        cosine[986] = 11'sd995;
        cosine[987] = 11'sd996;
        cosine[988] = 11'sd998;
        cosine[989] = 11'sd999;
        cosine[990] = 11'sd1000;
        cosine[991] = 11'sd1002;
        cosine[992] = 11'sd1003;
        cosine[993] = 11'sd1004;
        cosine[994] = 11'sd1005;
        cosine[995] = 11'sd1006;
        cosine[996] = 11'sd1007;
        cosine[997] = 11'sd1008;
        cosine[998] = 11'sd1010;
        cosine[999] = 11'sd1010;
        cosine[1000] = 11'sd1011;
        cosine[1001] = 11'sd1012;
        cosine[1002] = 11'sd1013;
        cosine[1003] = 11'sd1014;
        cosine[1004] = 11'sd1015;
        cosine[1005] = 11'sd1016;
        cosine[1006] = 11'sd1016;
        cosine[1007] = 11'sd1017;
        cosine[1008] = 11'sd1018;
        cosine[1009] = 11'sd1018;
        cosine[1010] = 11'sd1019;
        cosine[1011] = 11'sd1019;
        cosine[1012] = 11'sd1020;
        cosine[1013] = 11'sd1020;
        cosine[1014] = 11'sd1021;
        cosine[1015] = 11'sd1021;
        cosine[1016] = 11'sd1021;
        cosine[1017] = 11'sd1022;
        cosine[1018] = 11'sd1022;
        cosine[1019] = 11'sd1022;
        cosine[1020] = 11'sd1022;
        cosine[1021] = 11'sd1022;
        cosine[1022] = 11'sd1022;
        cosine[1023] = 11'sd1022;
    end

endmodule


