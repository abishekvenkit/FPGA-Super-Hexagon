module start_screen(input  logic Clk,
           input  logic [6:0] row_addr,
           output logic [159:0] columns);

    reg [159:0] img [0:119];

    always_ff @ (posedge Clk) begin
        columns <= img[row_addr];
    end

    initial begin
img[0] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[1] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[2] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[3] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[4] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[5] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[6] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[7] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[8] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[9] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[10] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[11] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[12] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[13] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[14] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[15] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[16] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[17] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[18] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[19] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[20] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[21] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[22] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[23] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[24] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[25] = 160'b0000000000000000000000000000000000000001111111111111110111111111111111100111111111111111001110000000001111001111111111111100000000000000000000000000000000000000;
img[26] = 160'b0000000000000000000000000000000000000011111111111111110111111111111111100111111111111111101111000000001111011111111111111110000000000000000000000000000000000000;
img[27] = 160'b0000000000000000000000000000000000000011111111111111110111111111111111100111111111111111101111000000001111011111111111111110000000000000000000000000000000000000;
img[28] = 160'b0000000000000000000000000000000000000011111111111111110111111111111111100111111111111111101111000000001111011111111111111110000000000000000000000000000000000000;
img[29] = 160'b0000000000000000000000000000000000000011110000000011110000000000000111100111000000000111101111000000001111000000000000001110000000000000000000000000000000000000;
img[30] = 160'b0000000000000000000000000000000000000011110000000011110000000000000111100111000000000111101111000000001111000000000000001110000000000000000000000000000000000000;
img[31] = 160'b0000000000000000000000000000000000000011110000000011110000000000000111100111000000000111101111000000001111000000000000011110000000000000000000000000000000000000;
img[32] = 160'b0000000000000000000000000000000000000011110000000011110111111111111111100111000000000111101111000000001111011111111111111110000000000000000000000000000000000000;
img[33] = 160'b0000000000000000000000000000000000000011110000000011110111111111111111100111100000000111101111000000001111011111111111111110000000000000000000000000000000000000;
img[34] = 160'b0000000000000000000000000000000000000011111111111111110111111111111111100111111111111111101111000000001111011111111111111110000000000000000000000000000000000000;
img[35] = 160'b0000000000000000000000000000000000000001111111111111110111111111111111100111111111111111101111000000001111011111111111111110000000000000000000000000000000000000;
img[36] = 160'b0000000000000000000000000000000000000011111111111111110000000000000111100111111111111111101111000000001111011110000000000000000000000000000000000000000000000000;
img[37] = 160'b0000000000000000000000000000000000000011111111111111110000000000000111100011111111111111101111000000001111011110000000000000000000000000000000000000000000000000;
img[38] = 160'b0000000000000000000000000000000000000011110000000011110111111111111111100000000000000111101111111111111111011111111111111110000000000000000000000000000000000000;
img[39] = 160'b0000000000000000000000000000000000000011110000000011110111111111111111100000000000000111101111111111111111011111111111111110000000000000000000000000000000000000;
img[40] = 160'b0000000000000000000000000000000000000011110000000011110111111111111111100000000000000111101111111111111111011111111111111110000000000000000000000000000000000000;
img[41] = 160'b0000000000000000000000000000000000000011110000000011110111111111111111000000000000000111101111111111111110001111111111111110000000000000000000000000000000000000;
img[42] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[43] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[44] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[45] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[46] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[47] = 160'b0000000000000000000001111111111111110011111111111111100111111111111111100111111111111111001110000000001111001111111111111110111100000000011100000000000000000000;
img[48] = 160'b0000000000000000000011111111111111110011111111111111110111111111111111100111111111111111001111000000001111011111111111111110111100000000011110000000000000000000;
img[49] = 160'b0000000000000000000011111111111111110011111111111111110111111111111111100111111111111111101111000000001111011111111111111110111100000000011110000000000000000000;
img[50] = 160'b0000000000000000000011111111111111110011111111111111110111111111111111100111111111111111101111000000001111011111111111111110111100000000011110000000000000000000;
img[51] = 160'b0000000000000000000011110000000001110011110000000011110000000000000111100111000000000111101111000000001111000000000000001110111100000000011110000000000000000000;
img[52] = 160'b0000000000000000000011110000000001110011110000000011110000000000000111100111000000000111101111000000001111000000000000001110111100000000011110000000000000000000;
img[53] = 160'b0000000000000000000011110000000001110011110000000011110000000000000111100111000000000111101111000000001111000000000000011110111110000000011110000000000000000000;
img[54] = 160'b0000000000000000000011110000000001110011110000000011110111100000000111100111000000000111101111111111111111011111111111111110111111111111111110000000000000000000;
img[55] = 160'b0000000000000000000011110000000001110011110000000011110111100000000111100111100000000111100111111111111110011111111111111110111111111111111110000000000000000000;
img[56] = 160'b0000000000000000000011110000000001110011110000000011110111100000000111100111111111111111101111111111111110011111111111111110111111111111111110000000000000000000;
img[57] = 160'b0000000000000000000011110000000001110011110000000011110111100000000111100111111111111111101111111111111111001111111111111110111111111111111110000000000000000000;
img[58] = 160'b0000000000000000000011110000000001110011110000000011110111100000000111100111111111111111101111000000001111000000000000001110111100000000011110000000000000000000;
img[59] = 160'b0000000000000000000011110000000001110011110000000011110111100000000111100111111111111111101111000000001111000000000000001110111100000000011110000000000000000000;
img[60] = 160'b0000000000000000000011110000000001110011111111111111110111111111111111100111000000000111101111000000001111011111111111111110111100000000011110000000000000000000;
img[61] = 160'b0000000000000000000011110000000001110011111111111111110111111111111111100111000000000111101111000000001111011111111111111110111100000000011110000000000000000000;
img[62] = 160'b0000000000000000000011110000000001110011111111111111110111111111111111100111000000000111101111000000001111011111111111111110111100000000011110000000000000000000;
img[63] = 160'b0000000000000000000011110000000001110001111111111111110011111111111111100111000000000111101111000000001111011111111111111100011100000000011110000000000000000000;
img[64] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[65] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[66] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[67] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[68] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[69] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[70] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[71] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[72] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[73] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[74] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[75] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[76] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[77] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[78] = 160'b0000000000000000000111111000000000001111100111110000000000000000001111100000000000000000001100000000000001111100011111001111110011111100111111000000000000000000;
img[79] = 160'b0000000000000000000011000000000000011001101100011000000000000000001100110000000000000000001110000000000011000110110011100000110110001101100011000000000000000000;
img[80] = 160'b0000000000000000000001100000000000011001101100011000000000000000001110000000000000000000001100000000000000000110000011100000110110001101100011000000000000000000;
img[81] = 160'b0000000000000000000011110000000000011101101100011000000000000000000111000000000000000000001100000000000001111100011111001111110111001101100011000000000000000000;
img[82] = 160'b0000000000000000000110000000000000001111101100011000000000000000000111100000000000000000001100000000000011000000110000000000110001111100111111000000000000000000;
img[83] = 160'b0000000000000000000110001100000000001101101100011000000000000110000001110000000000001100001100000000000011000110110011100000110011101100000011000000000000000000;
img[84] = 160'b0000000000000000000011111000000000011101100111110000000000000110001111110000000000001100011111000000000001111100011111001111110111001100000011000000000000000000;
img[85] = 160'b0000000000000000000000000000000000000000000000000000000000000011000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000;
img[86] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[87] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[88] = 160'b0000000000000000000000000000000000000000000000000111111100111110001111100011111001100011001110000000000001111100111111000000000000000000000000000000000000000000;
img[89] = 160'b0000000000000000000000000000000000000000000000000000001101100111011000110110001101100011011011000000000011000110001100000000000000000000000000000000000000000000;
img[90] = 160'b0000000000000000000000000000000000000000000000000000001100000111011000110110001101100011000001100000000011000110001100000000000000000000000000000000000000000000;
img[91] = 160'b0000000000000000000000000000000000000000000000000011111100111110011000110110001101111111000001100000000011000110001100000000000000000000000000000000000000000000;
img[92] = 160'b0000000000000000000000000000000000000000000000000000001101100000011000110110001101100011000001100000000011000110001100000000000000000000000000000000000000000000;
img[93] = 160'b0000000000000000000000000000000000000000000000000000001101100111011000110110001101100011011011000000000011000110001100000000000000000000000000000000000000000000;
img[94] = 160'b0000000000000000000000000000000000000000000000000111111100111110001111100011111001100011001110000000000001111100001100000000000000000000000000000000000000000000;
img[95] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[96] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[97] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[98] = 160'b0000000000000000000000000000000000000000001100110011111100000011001100110011110001111110011111101111111011111100001111100000000000000000000000000000000000000000;
img[99] = 160'b0000000000000000000000000000000000000000001100110000110000000011001100110110011000011000000001100000011000110000011001100000000000000000000000000000000000000000;
img[100] = 160'b0000000000000000000000000000000000000000001100110000110000000011001100110000001100011000000001100000011000110000110001100000000000000000000000000000000000000000;
img[101] = 160'b0000000000000000000000000000000000000000000111100000110000000011001100110000001100011000001111100111111000110000110001100000000000000000000000000000000000000000;
img[102] = 160'b0000000000000000000000000000000000000000000011000000110000000011001100110000001100011000000001100000011000110000110001100000000000000000000000000000000000000000;
img[103] = 160'b0000000000000000000000000000000000000000000011000000110000000011001100110110011000011000000001100000011000110000011001100000000000000000000000000000000000000000;
img[104] = 160'b0000000000000000000000000000000000000000000011000000110000111111000111100011110001111110000001100000011011111100001111100000000000000000000000000000000000000000;
img[105] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[106] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[107] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[108] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[109] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[110] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[111] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[112] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[113] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[114] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[115] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[116] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[117] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[118] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
img[119] = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
endmodule