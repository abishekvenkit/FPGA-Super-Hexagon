module sin (input  logic        Clk,
            input  logic  [9:0] angle,
            output logic [20:0] answer);
    
    reg signed [10:0] sine [0:1023];
    logic signed [10:0] answer_10;

    assign answer = {{10{answer_10[10]}}, answer_10};
    always_ff @ (posedge Clk) begin
        answer_10 <= sine[angle];
    end

    initial begin
        sine[0] = 11'sd0;
        sine[1] = 11'sd6;
        sine[2] = 11'sd12;
        sine[3] = 11'sd18;
        sine[4] = 11'sd25;
        sine[5] = 11'sd31;
        sine[6] = 11'sd37;
        sine[7] = 11'sd43;
        sine[8] = 11'sd50;
        sine[9] = 11'sd56;
        sine[10] = 11'sd62;
        sine[11] = 11'sd68;
        sine[12] = 11'sd75;
        sine[13] = 11'sd81;
        sine[14] = 11'sd87;
        sine[15] = 11'sd94;
        sine[16] = 11'sd100;
        sine[17] = 11'sd106;
        sine[18] = 11'sd112;
        sine[19] = 11'sd118;
        sine[20] = 11'sd125;
        sine[21] = 11'sd131;
        sine[22] = 11'sd137;
        sine[23] = 11'sd143;
        sine[24] = 11'sd150;
        sine[25] = 11'sd156;
        sine[26] = 11'sd162;
        sine[27] = 11'sd168;
        sine[28] = 11'sd174;
        sine[29] = 11'sd181;
        sine[30] = 11'sd187;
        sine[31] = 11'sd193;
        sine[32] = 11'sd199;
        sine[33] = 11'sd205;
        sine[34] = 11'sd211;
        sine[35] = 11'sd218;
        sine[36] = 11'sd224;
        sine[37] = 11'sd230;
        sine[38] = 11'sd236;
        sine[39] = 11'sd242;
        sine[40] = 11'sd248;
        sine[41] = 11'sd254;
        sine[42] = 11'sd260;
        sine[43] = 11'sd266;
        sine[44] = 11'sd272;
        sine[45] = 11'sd278;
        sine[46] = 11'sd284;
        sine[47] = 11'sd290;
        sine[48] = 11'sd296;
        sine[49] = 11'sd302;
        sine[50] = 11'sd308;
        sine[51] = 11'sd314;
        sine[52] = 11'sd320;
        sine[53] = 11'sd326;
        sine[54] = 11'sd332;
        sine[55] = 11'sd338;
        sine[56] = 11'sd344;
        sine[57] = 11'sd350;
        sine[58] = 11'sd356;
        sine[59] = 11'sd362;
        sine[60] = 11'sd368;
        sine[61] = 11'sd374;
        sine[62] = 11'sd379;
        sine[63] = 11'sd385;
        sine[64] = 11'sd391;
        sine[65] = 11'sd397;
        sine[66] = 11'sd403;
        sine[67] = 11'sd408;
        sine[68] = 11'sd414;
        sine[69] = 11'sd420;
        sine[70] = 11'sd426;
        sine[71] = 11'sd431;
        sine[72] = 11'sd437;
        sine[73] = 11'sd443;
        sine[74] = 11'sd448;
        sine[75] = 11'sd454;
        sine[76] = 11'sd459;
        sine[77] = 11'sd465;
        sine[78] = 11'sd471;
        sine[79] = 11'sd476;
        sine[80] = 11'sd482;
        sine[81] = 11'sd487;
        sine[82] = 11'sd493;
        sine[83] = 11'sd498;
        sine[84] = 11'sd504;
        sine[85] = 11'sd509;
        sine[86] = 11'sd515;
        sine[87] = 11'sd520;
        sine[88] = 11'sd525;
        sine[89] = 11'sd531;
        sine[90] = 11'sd536;
        sine[91] = 11'sd541;
        sine[92] = 11'sd547;
        sine[93] = 11'sd552;
        sine[94] = 11'sd557;
        sine[95] = 11'sd563;
        sine[96] = 11'sd568;
        sine[97] = 11'sd573;
        sine[98] = 11'sd578;
        sine[99] = 11'sd583;
        sine[100] = 11'sd589;
        sine[101] = 11'sd594;
        sine[102] = 11'sd599;
        sine[103] = 11'sd604;
        sine[104] = 11'sd609;
        sine[105] = 11'sd614;
        sine[106] = 11'sd619;
        sine[107] = 11'sd624;
        sine[108] = 11'sd629;
        sine[109] = 11'sd634;
        sine[110] = 11'sd639;
        sine[111] = 11'sd644;
        sine[112] = 11'sd648;
        sine[113] = 11'sd653;
        sine[114] = 11'sd658;
        sine[115] = 11'sd663;
        sine[116] = 11'sd668;
        sine[117] = 11'sd672;
        sine[118] = 11'sd677;
        sine[119] = 11'sd682;
        sine[120] = 11'sd687;
        sine[121] = 11'sd691;
        sine[122] = 11'sd696;
        sine[123] = 11'sd700;
        sine[124] = 11'sd705;
        sine[125] = 11'sd709;
        sine[126] = 11'sd714;
        sine[127] = 11'sd718;
        sine[128] = 11'sd723;
        sine[129] = 11'sd727;
        sine[130] = 11'sd732;
        sine[131] = 11'sd736;
        sine[132] = 11'sd740;
        sine[133] = 11'sd745;
        sine[134] = 11'sd749;
        sine[135] = 11'sd753;
        sine[136] = 11'sd757;
        sine[137] = 11'sd762;
        sine[138] = 11'sd766;
        sine[139] = 11'sd770;
        sine[140] = 11'sd774;
        sine[141] = 11'sd778;
        sine[142] = 11'sd782;
        sine[143] = 11'sd786;
        sine[144] = 11'sd790;
        sine[145] = 11'sd794;
        sine[146] = 11'sd798;
        sine[147] = 11'sd802;
        sine[148] = 11'sd806;
        sine[149] = 11'sd810;
        sine[150] = 11'sd814;
        sine[151] = 11'sd817;
        sine[152] = 11'sd821;
        sine[153] = 11'sd825;
        sine[154] = 11'sd829;
        sine[155] = 11'sd832;
        sine[156] = 11'sd836;
        sine[157] = 11'sd839;
        sine[158] = 11'sd843;
        sine[159] = 11'sd847;
        sine[160] = 11'sd850;
        sine[161] = 11'sd854;
        sine[162] = 11'sd857;
        sine[163] = 11'sd860;
        sine[164] = 11'sd864;
        sine[165] = 11'sd867;
        sine[166] = 11'sd870;
        sine[167] = 11'sd874;
        sine[168] = 11'sd877;
        sine[169] = 11'sd880;
        sine[170] = 11'sd883;
        sine[171] = 11'sd886;
        sine[172] = 11'sd890;
        sine[173] = 11'sd893;
        sine[174] = 11'sd896;
        sine[175] = 11'sd899;
        sine[176] = 11'sd902;
        sine[177] = 11'sd905;
        sine[178] = 11'sd908;
        sine[179] = 11'sd910;
        sine[180] = 11'sd913;
        sine[181] = 11'sd916;
        sine[182] = 11'sd919;
        sine[183] = 11'sd922;
        sine[184] = 11'sd924;
        sine[185] = 11'sd927;
        sine[186] = 11'sd930;
        sine[187] = 11'sd932;
        sine[188] = 11'sd935;
        sine[189] = 11'sd937;
        sine[190] = 11'sd940;
        sine[191] = 11'sd942;
        sine[192] = 11'sd945;
        sine[193] = 11'sd947;
        sine[194] = 11'sd949;
        sine[195] = 11'sd952;
        sine[196] = 11'sd954;
        sine[197] = 11'sd956;
        sine[198] = 11'sd958;
        sine[199] = 11'sd961;
        sine[200] = 11'sd963;
        sine[201] = 11'sd965;
        sine[202] = 11'sd967;
        sine[203] = 11'sd969;
        sine[204] = 11'sd971;
        sine[205] = 11'sd973;
        sine[206] = 11'sd975;
        sine[207] = 11'sd977;
        sine[208] = 11'sd978;
        sine[209] = 11'sd980;
        sine[210] = 11'sd982;
        sine[211] = 11'sd984;
        sine[212] = 11'sd985;
        sine[213] = 11'sd987;
        sine[214] = 11'sd989;
        sine[215] = 11'sd990;
        sine[216] = 11'sd992;
        sine[217] = 11'sd993;
        sine[218] = 11'sd995;
        sine[219] = 11'sd996;
        sine[220] = 11'sd998;
        sine[221] = 11'sd999;
        sine[222] = 11'sd1000;
        sine[223] = 11'sd1002;
        sine[224] = 11'sd1003;
        sine[225] = 11'sd1004;
        sine[226] = 11'sd1005;
        sine[227] = 11'sd1006;
        sine[228] = 11'sd1007;
        sine[229] = 11'sd1008;
        sine[230] = 11'sd1010;
        sine[231] = 11'sd1010;
        sine[232] = 11'sd1011;
        sine[233] = 11'sd1012;
        sine[234] = 11'sd1013;
        sine[235] = 11'sd1014;
        sine[236] = 11'sd1015;
        sine[237] = 11'sd1016;
        sine[238] = 11'sd1016;
        sine[239] = 11'sd1017;
        sine[240] = 11'sd1018;
        sine[241] = 11'sd1018;
        sine[242] = 11'sd1019;
        sine[243] = 11'sd1019;
        sine[244] = 11'sd1020;
        sine[245] = 11'sd1020;
        sine[246] = 11'sd1021;
        sine[247] = 11'sd1021;
        sine[248] = 11'sd1021;
        sine[249] = 11'sd1022;
        sine[250] = 11'sd1022;
        sine[251] = 11'sd1022;
        sine[252] = 11'sd1022;
        sine[253] = 11'sd1022;
        sine[254] = 11'sd1022;
        sine[255] = 11'sd1022;
        sine[256] = 11'sd1023;
        sine[257] = 11'sd1022;
        sine[258] = 11'sd1022;
        sine[259] = 11'sd1022;
        sine[260] = 11'sd1022;
        sine[261] = 11'sd1022;
        sine[262] = 11'sd1022;
        sine[263] = 11'sd1022;
        sine[264] = 11'sd1021;
        sine[265] = 11'sd1021;
        sine[266] = 11'sd1021;
        sine[267] = 11'sd1020;
        sine[268] = 11'sd1020;
        sine[269] = 11'sd1019;
        sine[270] = 11'sd1019;
        sine[271] = 11'sd1018;
        sine[272] = 11'sd1018;
        sine[273] = 11'sd1017;
        sine[274] = 11'sd1016;
        sine[275] = 11'sd1016;
        sine[276] = 11'sd1015;
        sine[277] = 11'sd1014;
        sine[278] = 11'sd1013;
        sine[279] = 11'sd1012;
        sine[280] = 11'sd1011;
        sine[281] = 11'sd1010;
        sine[282] = 11'sd1010;
        sine[283] = 11'sd1008;
        sine[284] = 11'sd1007;
        sine[285] = 11'sd1006;
        sine[286] = 11'sd1005;
        sine[287] = 11'sd1004;
        sine[288] = 11'sd1003;
        sine[289] = 11'sd1002;
        sine[290] = 11'sd1000;
        sine[291] = 11'sd999;
        sine[292] = 11'sd998;
        sine[293] = 11'sd996;
        sine[294] = 11'sd995;
        sine[295] = 11'sd993;
        sine[296] = 11'sd992;
        sine[297] = 11'sd990;
        sine[298] = 11'sd989;
        sine[299] = 11'sd987;
        sine[300] = 11'sd985;
        sine[301] = 11'sd984;
        sine[302] = 11'sd982;
        sine[303] = 11'sd980;
        sine[304] = 11'sd978;
        sine[305] = 11'sd977;
        sine[306] = 11'sd975;
        sine[307] = 11'sd973;
        sine[308] = 11'sd971;
        sine[309] = 11'sd969;
        sine[310] = 11'sd967;
        sine[311] = 11'sd965;
        sine[312] = 11'sd963;
        sine[313] = 11'sd961;
        sine[314] = 11'sd958;
        sine[315] = 11'sd956;
        sine[316] = 11'sd954;
        sine[317] = 11'sd952;
        sine[318] = 11'sd949;
        sine[319] = 11'sd947;
        sine[320] = 11'sd945;
        sine[321] = 11'sd942;
        sine[322] = 11'sd940;
        sine[323] = 11'sd937;
        sine[324] = 11'sd935;
        sine[325] = 11'sd932;
        sine[326] = 11'sd930;
        sine[327] = 11'sd927;
        sine[328] = 11'sd924;
        sine[329] = 11'sd922;
        sine[330] = 11'sd919;
        sine[331] = 11'sd916;
        sine[332] = 11'sd913;
        sine[333] = 11'sd910;
        sine[334] = 11'sd908;
        sine[335] = 11'sd905;
        sine[336] = 11'sd902;
        sine[337] = 11'sd899;
        sine[338] = 11'sd896;
        sine[339] = 11'sd893;
        sine[340] = 11'sd890;
        sine[341] = 11'sd886;
        sine[342] = 11'sd883;
        sine[343] = 11'sd880;
        sine[344] = 11'sd877;
        sine[345] = 11'sd874;
        sine[346] = 11'sd870;
        sine[347] = 11'sd867;
        sine[348] = 11'sd864;
        sine[349] = 11'sd860;
        sine[350] = 11'sd857;
        sine[351] = 11'sd854;
        sine[352] = 11'sd850;
        sine[353] = 11'sd847;
        sine[354] = 11'sd843;
        sine[355] = 11'sd839;
        sine[356] = 11'sd836;
        sine[357] = 11'sd832;
        sine[358] = 11'sd829;
        sine[359] = 11'sd825;
        sine[360] = 11'sd821;
        sine[361] = 11'sd817;
        sine[362] = 11'sd814;
        sine[363] = 11'sd810;
        sine[364] = 11'sd806;
        sine[365] = 11'sd802;
        sine[366] = 11'sd798;
        sine[367] = 11'sd794;
        sine[368] = 11'sd790;
        sine[369] = 11'sd786;
        sine[370] = 11'sd782;
        sine[371] = 11'sd778;
        sine[372] = 11'sd774;
        sine[373] = 11'sd770;
        sine[374] = 11'sd766;
        sine[375] = 11'sd762;
        sine[376] = 11'sd757;
        sine[377] = 11'sd753;
        sine[378] = 11'sd749;
        sine[379] = 11'sd745;
        sine[380] = 11'sd740;
        sine[381] = 11'sd736;
        sine[382] = 11'sd732;
        sine[383] = 11'sd727;
        sine[384] = 11'sd723;
        sine[385] = 11'sd718;
        sine[386] = 11'sd714;
        sine[387] = 11'sd709;
        sine[388] = 11'sd705;
        sine[389] = 11'sd700;
        sine[390] = 11'sd696;
        sine[391] = 11'sd691;
        sine[392] = 11'sd687;
        sine[393] = 11'sd682;
        sine[394] = 11'sd677;
        sine[395] = 11'sd672;
        sine[396] = 11'sd668;
        sine[397] = 11'sd663;
        sine[398] = 11'sd658;
        sine[399] = 11'sd653;
        sine[400] = 11'sd648;
        sine[401] = 11'sd644;
        sine[402] = 11'sd639;
        sine[403] = 11'sd634;
        sine[404] = 11'sd629;
        sine[405] = 11'sd624;
        sine[406] = 11'sd619;
        sine[407] = 11'sd614;
        sine[408] = 11'sd609;
        sine[409] = 11'sd604;
        sine[410] = 11'sd599;
        sine[411] = 11'sd594;
        sine[412] = 11'sd589;
        sine[413] = 11'sd583;
        sine[414] = 11'sd578;
        sine[415] = 11'sd573;
        sine[416] = 11'sd568;
        sine[417] = 11'sd563;
        sine[418] = 11'sd557;
        sine[419] = 11'sd552;
        sine[420] = 11'sd547;
        sine[421] = 11'sd541;
        sine[422] = 11'sd536;
        sine[423] = 11'sd531;
        sine[424] = 11'sd525;
        sine[425] = 11'sd520;
        sine[426] = 11'sd515;
        sine[427] = 11'sd509;
        sine[428] = 11'sd504;
        sine[429] = 11'sd498;
        sine[430] = 11'sd493;
        sine[431] = 11'sd487;
        sine[432] = 11'sd482;
        sine[433] = 11'sd476;
        sine[434] = 11'sd471;
        sine[435] = 11'sd465;
        sine[436] = 11'sd459;
        sine[437] = 11'sd454;
        sine[438] = 11'sd448;
        sine[439] = 11'sd443;
        sine[440] = 11'sd437;
        sine[441] = 11'sd431;
        sine[442] = 11'sd426;
        sine[443] = 11'sd420;
        sine[444] = 11'sd414;
        sine[445] = 11'sd408;
        sine[446] = 11'sd403;
        sine[447] = 11'sd397;
        sine[448] = 11'sd391;
        sine[449] = 11'sd385;
        sine[450] = 11'sd379;
        sine[451] = 11'sd374;
        sine[452] = 11'sd368;
        sine[453] = 11'sd362;
        sine[454] = 11'sd356;
        sine[455] = 11'sd350;
        sine[456] = 11'sd344;
        sine[457] = 11'sd338;
        sine[458] = 11'sd332;
        sine[459] = 11'sd326;
        sine[460] = 11'sd320;
        sine[461] = 11'sd314;
        sine[462] = 11'sd308;
        sine[463] = 11'sd302;
        sine[464] = 11'sd296;
        sine[465] = 11'sd290;
        sine[466] = 11'sd284;
        sine[467] = 11'sd278;
        sine[468] = 11'sd272;
        sine[469] = 11'sd266;
        sine[470] = 11'sd260;
        sine[471] = 11'sd254;
        sine[472] = 11'sd248;
        sine[473] = 11'sd242;
        sine[474] = 11'sd236;
        sine[475] = 11'sd230;
        sine[476] = 11'sd224;
        sine[477] = 11'sd218;
        sine[478] = 11'sd211;
        sine[479] = 11'sd205;
        sine[480] = 11'sd199;
        sine[481] = 11'sd193;
        sine[482] = 11'sd187;
        sine[483] = 11'sd181;
        sine[484] = 11'sd174;
        sine[485] = 11'sd168;
        sine[486] = 11'sd162;
        sine[487] = 11'sd156;
        sine[488] = 11'sd150;
        sine[489] = 11'sd143;
        sine[490] = 11'sd137;
        sine[491] = 11'sd131;
        sine[492] = 11'sd125;
        sine[493] = 11'sd118;
        sine[494] = 11'sd112;
        sine[495] = 11'sd106;
        sine[496] = 11'sd100;
        sine[497] = 11'sd94;
        sine[498] = 11'sd87;
        sine[499] = 11'sd81;
        sine[500] = 11'sd75;
        sine[501] = 11'sd68;
        sine[502] = 11'sd62;
        sine[503] = 11'sd56;
        sine[504] = 11'sd50;
        sine[505] = 11'sd43;
        sine[506] = 11'sd37;
        sine[507] = 11'sd31;
        sine[508] = 11'sd25;
        sine[509] = 11'sd18;
        sine[510] = 11'sd12;
        sine[511] = 11'sd6;
        sine[512] = 11'sd0;
        sine[513] = -11'sd6;
        sine[514] = -11'sd12;
        sine[515] = -11'sd18;
        sine[516] = -11'sd25;
        sine[517] = -11'sd31;
        sine[518] = -11'sd37;
        sine[519] = -11'sd43;
        sine[520] = -11'sd50;
        sine[521] = -11'sd56;
        sine[522] = -11'sd62;
        sine[523] = -11'sd68;
        sine[524] = -11'sd75;
        sine[525] = -11'sd81;
        sine[526] = -11'sd87;
        sine[527] = -11'sd94;
        sine[528] = -11'sd100;
        sine[529] = -11'sd106;
        sine[530] = -11'sd112;
        sine[531] = -11'sd118;
        sine[532] = -11'sd125;
        sine[533] = -11'sd131;
        sine[534] = -11'sd137;
        sine[535] = -11'sd143;
        sine[536] = -11'sd150;
        sine[537] = -11'sd156;
        sine[538] = -11'sd162;
        sine[539] = -11'sd168;
        sine[540] = -11'sd174;
        sine[541] = -11'sd181;
        sine[542] = -11'sd187;
        sine[543] = -11'sd193;
        sine[544] = -11'sd199;
        sine[545] = -11'sd205;
        sine[546] = -11'sd211;
        sine[547] = -11'sd218;
        sine[548] = -11'sd224;
        sine[549] = -11'sd230;
        sine[550] = -11'sd236;
        sine[551] = -11'sd242;
        sine[552] = -11'sd248;
        sine[553] = -11'sd254;
        sine[554] = -11'sd260;
        sine[555] = -11'sd266;
        sine[556] = -11'sd272;
        sine[557] = -11'sd278;
        sine[558] = -11'sd284;
        sine[559] = -11'sd290;
        sine[560] = -11'sd296;
        sine[561] = -11'sd302;
        sine[562] = -11'sd308;
        sine[563] = -11'sd314;
        sine[564] = -11'sd320;
        sine[565] = -11'sd326;
        sine[566] = -11'sd332;
        sine[567] = -11'sd338;
        sine[568] = -11'sd344;
        sine[569] = -11'sd350;
        sine[570] = -11'sd356;
        sine[571] = -11'sd362;
        sine[572] = -11'sd368;
        sine[573] = -11'sd374;
        sine[574] = -11'sd379;
        sine[575] = -11'sd385;
        sine[576] = -11'sd391;
        sine[577] = -11'sd397;
        sine[578] = -11'sd403;
        sine[579] = -11'sd408;
        sine[580] = -11'sd414;
        sine[581] = -11'sd420;
        sine[582] = -11'sd426;
        sine[583] = -11'sd431;
        sine[584] = -11'sd437;
        sine[585] = -11'sd443;
        sine[586] = -11'sd448;
        sine[587] = -11'sd454;
        sine[588] = -11'sd459;
        sine[589] = -11'sd465;
        sine[590] = -11'sd471;
        sine[591] = -11'sd476;
        sine[592] = -11'sd482;
        sine[593] = -11'sd487;
        sine[594] = -11'sd493;
        sine[595] = -11'sd498;
        sine[596] = -11'sd504;
        sine[597] = -11'sd509;
        sine[598] = -11'sd515;
        sine[599] = -11'sd520;
        sine[600] = -11'sd525;
        sine[601] = -11'sd531;
        sine[602] = -11'sd536;
        sine[603] = -11'sd541;
        sine[604] = -11'sd547;
        sine[605] = -11'sd552;
        sine[606] = -11'sd557;
        sine[607] = -11'sd563;
        sine[608] = -11'sd568;
        sine[609] = -11'sd573;
        sine[610] = -11'sd578;
        sine[611] = -11'sd583;
        sine[612] = -11'sd589;
        sine[613] = -11'sd594;
        sine[614] = -11'sd599;
        sine[615] = -11'sd604;
        sine[616] = -11'sd609;
        sine[617] = -11'sd614;
        sine[618] = -11'sd619;
        sine[619] = -11'sd624;
        sine[620] = -11'sd629;
        sine[621] = -11'sd634;
        sine[622] = -11'sd639;
        sine[623] = -11'sd644;
        sine[624] = -11'sd648;
        sine[625] = -11'sd653;
        sine[626] = -11'sd658;
        sine[627] = -11'sd663;
        sine[628] = -11'sd668;
        sine[629] = -11'sd672;
        sine[630] = -11'sd677;
        sine[631] = -11'sd682;
        sine[632] = -11'sd687;
        sine[633] = -11'sd691;
        sine[634] = -11'sd696;
        sine[635] = -11'sd700;
        sine[636] = -11'sd705;
        sine[637] = -11'sd709;
        sine[638] = -11'sd714;
        sine[639] = -11'sd718;
        sine[640] = -11'sd723;
        sine[641] = -11'sd727;
        sine[642] = -11'sd732;
        sine[643] = -11'sd736;
        sine[644] = -11'sd740;
        sine[645] = -11'sd745;
        sine[646] = -11'sd749;
        sine[647] = -11'sd753;
        sine[648] = -11'sd757;
        sine[649] = -11'sd762;
        sine[650] = -11'sd766;
        sine[651] = -11'sd770;
        sine[652] = -11'sd774;
        sine[653] = -11'sd778;
        sine[654] = -11'sd782;
        sine[655] = -11'sd786;
        sine[656] = -11'sd790;
        sine[657] = -11'sd794;
        sine[658] = -11'sd798;
        sine[659] = -11'sd802;
        sine[660] = -11'sd806;
        sine[661] = -11'sd810;
        sine[662] = -11'sd814;
        sine[663] = -11'sd817;
        sine[664] = -11'sd821;
        sine[665] = -11'sd825;
        sine[666] = -11'sd829;
        sine[667] = -11'sd832;
        sine[668] = -11'sd836;
        sine[669] = -11'sd839;
        sine[670] = -11'sd843;
        sine[671] = -11'sd847;
        sine[672] = -11'sd850;
        sine[673] = -11'sd854;
        sine[674] = -11'sd857;
        sine[675] = -11'sd860;
        sine[676] = -11'sd864;
        sine[677] = -11'sd867;
        sine[678] = -11'sd870;
        sine[679] = -11'sd874;
        sine[680] = -11'sd877;
        sine[681] = -11'sd880;
        sine[682] = -11'sd883;
        sine[683] = -11'sd886;
        sine[684] = -11'sd890;
        sine[685] = -11'sd893;
        sine[686] = -11'sd896;
        sine[687] = -11'sd899;
        sine[688] = -11'sd902;
        sine[689] = -11'sd905;
        sine[690] = -11'sd908;
        sine[691] = -11'sd910;
        sine[692] = -11'sd913;
        sine[693] = -11'sd916;
        sine[694] = -11'sd919;
        sine[695] = -11'sd922;
        sine[696] = -11'sd924;
        sine[697] = -11'sd927;
        sine[698] = -11'sd930;
        sine[699] = -11'sd932;
        sine[700] = -11'sd935;
        sine[701] = -11'sd937;
        sine[702] = -11'sd940;
        sine[703] = -11'sd942;
        sine[704] = -11'sd945;
        sine[705] = -11'sd947;
        sine[706] = -11'sd949;
        sine[707] = -11'sd952;
        sine[708] = -11'sd954;
        sine[709] = -11'sd956;
        sine[710] = -11'sd958;
        sine[711] = -11'sd961;
        sine[712] = -11'sd963;
        sine[713] = -11'sd965;
        sine[714] = -11'sd967;
        sine[715] = -11'sd969;
        sine[716] = -11'sd971;
        sine[717] = -11'sd973;
        sine[718] = -11'sd975;
        sine[719] = -11'sd977;
        sine[720] = -11'sd978;
        sine[721] = -11'sd980;
        sine[722] = -11'sd982;
        sine[723] = -11'sd984;
        sine[724] = -11'sd985;
        sine[725] = -11'sd987;
        sine[726] = -11'sd989;
        sine[727] = -11'sd990;
        sine[728] = -11'sd992;
        sine[729] = -11'sd993;
        sine[730] = -11'sd995;
        sine[731] = -11'sd996;
        sine[732] = -11'sd998;
        sine[733] = -11'sd999;
        sine[734] = -11'sd1000;
        sine[735] = -11'sd1002;
        sine[736] = -11'sd1003;
        sine[737] = -11'sd1004;
        sine[738] = -11'sd1005;
        sine[739] = -11'sd1006;
        sine[740] = -11'sd1007;
        sine[741] = -11'sd1008;
        sine[742] = -11'sd1010;
        sine[743] = -11'sd1010;
        sine[744] = -11'sd1011;
        sine[745] = -11'sd1012;
        sine[746] = -11'sd1013;
        sine[747] = -11'sd1014;
        sine[748] = -11'sd1015;
        sine[749] = -11'sd1016;
        sine[750] = -11'sd1016;
        sine[751] = -11'sd1017;
        sine[752] = -11'sd1018;
        sine[753] = -11'sd1018;
        sine[754] = -11'sd1019;
        sine[755] = -11'sd1019;
        sine[756] = -11'sd1020;
        sine[757] = -11'sd1020;
        sine[758] = -11'sd1021;
        sine[759] = -11'sd1021;
        sine[760] = -11'sd1021;
        sine[761] = -11'sd1022;
        sine[762] = -11'sd1022;
        sine[763] = -11'sd1022;
        sine[764] = -11'sd1022;
        sine[765] = -11'sd1022;
        sine[766] = -11'sd1022;
        sine[767] = -11'sd1022;
        sine[768] = -11'sd1023;
        sine[769] = -11'sd1022;
        sine[770] = -11'sd1022;
        sine[771] = -11'sd1022;
        sine[772] = -11'sd1022;
        sine[773] = -11'sd1022;
        sine[774] = -11'sd1022;
        sine[775] = -11'sd1022;
        sine[776] = -11'sd1021;
        sine[777] = -11'sd1021;
        sine[778] = -11'sd1021;
        sine[779] = -11'sd1020;
        sine[780] = -11'sd1020;
        sine[781] = -11'sd1019;
        sine[782] = -11'sd1019;
        sine[783] = -11'sd1018;
        sine[784] = -11'sd1018;
        sine[785] = -11'sd1017;
        sine[786] = -11'sd1016;
        sine[787] = -11'sd1016;
        sine[788] = -11'sd1015;
        sine[789] = -11'sd1014;
        sine[790] = -11'sd1013;
        sine[791] = -11'sd1012;
        sine[792] = -11'sd1011;
        sine[793] = -11'sd1010;
        sine[794] = -11'sd1010;
        sine[795] = -11'sd1008;
        sine[796] = -11'sd1007;
        sine[797] = -11'sd1006;
        sine[798] = -11'sd1005;
        sine[799] = -11'sd1004;
        sine[800] = -11'sd1003;
        sine[801] = -11'sd1002;
        sine[802] = -11'sd1000;
        sine[803] = -11'sd999;
        sine[804] = -11'sd998;
        sine[805] = -11'sd996;
        sine[806] = -11'sd995;
        sine[807] = -11'sd993;
        sine[808] = -11'sd992;
        sine[809] = -11'sd990;
        sine[810] = -11'sd989;
        sine[811] = -11'sd987;
        sine[812] = -11'sd985;
        sine[813] = -11'sd984;
        sine[814] = -11'sd982;
        sine[815] = -11'sd980;
        sine[816] = -11'sd978;
        sine[817] = -11'sd977;
        sine[818] = -11'sd975;
        sine[819] = -11'sd973;
        sine[820] = -11'sd971;
        sine[821] = -11'sd969;
        sine[822] = -11'sd967;
        sine[823] = -11'sd965;
        sine[824] = -11'sd963;
        sine[825] = -11'sd961;
        sine[826] = -11'sd958;
        sine[827] = -11'sd956;
        sine[828] = -11'sd954;
        sine[829] = -11'sd952;
        sine[830] = -11'sd949;
        sine[831] = -11'sd947;
        sine[832] = -11'sd945;
        sine[833] = -11'sd942;
        sine[834] = -11'sd940;
        sine[835] = -11'sd937;
        sine[836] = -11'sd935;
        sine[837] = -11'sd932;
        sine[838] = -11'sd930;
        sine[839] = -11'sd927;
        sine[840] = -11'sd924;
        sine[841] = -11'sd922;
        sine[842] = -11'sd919;
        sine[843] = -11'sd916;
        sine[844] = -11'sd913;
        sine[845] = -11'sd910;
        sine[846] = -11'sd908;
        sine[847] = -11'sd905;
        sine[848] = -11'sd902;
        sine[849] = -11'sd899;
        sine[850] = -11'sd896;
        sine[851] = -11'sd893;
        sine[852] = -11'sd890;
        sine[853] = -11'sd886;
        sine[854] = -11'sd883;
        sine[855] = -11'sd880;
        sine[856] = -11'sd877;
        sine[857] = -11'sd874;
        sine[858] = -11'sd870;
        sine[859] = -11'sd867;
        sine[860] = -11'sd864;
        sine[861] = -11'sd860;
        sine[862] = -11'sd857;
        sine[863] = -11'sd854;
        sine[864] = -11'sd850;
        sine[865] = -11'sd847;
        sine[866] = -11'sd843;
        sine[867] = -11'sd839;
        sine[868] = -11'sd836;
        sine[869] = -11'sd832;
        sine[870] = -11'sd829;
        sine[871] = -11'sd825;
        sine[872] = -11'sd821;
        sine[873] = -11'sd817;
        sine[874] = -11'sd814;
        sine[875] = -11'sd810;
        sine[876] = -11'sd806;
        sine[877] = -11'sd802;
        sine[878] = -11'sd798;
        sine[879] = -11'sd794;
        sine[880] = -11'sd790;
        sine[881] = -11'sd786;
        sine[882] = -11'sd782;
        sine[883] = -11'sd778;
        sine[884] = -11'sd774;
        sine[885] = -11'sd770;
        sine[886] = -11'sd766;
        sine[887] = -11'sd762;
        sine[888] = -11'sd757;
        sine[889] = -11'sd753;
        sine[890] = -11'sd749;
        sine[891] = -11'sd745;
        sine[892] = -11'sd740;
        sine[893] = -11'sd736;
        sine[894] = -11'sd732;
        sine[895] = -11'sd727;
        sine[896] = -11'sd723;
        sine[897] = -11'sd718;
        sine[898] = -11'sd714;
        sine[899] = -11'sd709;
        sine[900] = -11'sd705;
        sine[901] = -11'sd700;
        sine[902] = -11'sd696;
        sine[903] = -11'sd691;
        sine[904] = -11'sd687;
        sine[905] = -11'sd682;
        sine[906] = -11'sd677;
        sine[907] = -11'sd672;
        sine[908] = -11'sd668;
        sine[909] = -11'sd663;
        sine[910] = -11'sd658;
        sine[911] = -11'sd653;
        sine[912] = -11'sd648;
        sine[913] = -11'sd644;
        sine[914] = -11'sd639;
        sine[915] = -11'sd634;
        sine[916] = -11'sd629;
        sine[917] = -11'sd624;
        sine[918] = -11'sd619;
        sine[919] = -11'sd614;
        sine[920] = -11'sd609;
        sine[921] = -11'sd604;
        sine[922] = -11'sd599;
        sine[923] = -11'sd594;
        sine[924] = -11'sd589;
        sine[925] = -11'sd583;
        sine[926] = -11'sd578;
        sine[927] = -11'sd573;
        sine[928] = -11'sd568;
        sine[929] = -11'sd563;
        sine[930] = -11'sd557;
        sine[931] = -11'sd552;
        sine[932] = -11'sd547;
        sine[933] = -11'sd541;
        sine[934] = -11'sd536;
        sine[935] = -11'sd531;
        sine[936] = -11'sd525;
        sine[937] = -11'sd520;
        sine[938] = -11'sd515;
        sine[939] = -11'sd509;
        sine[940] = -11'sd504;
        sine[941] = -11'sd498;
        sine[942] = -11'sd493;
        sine[943] = -11'sd487;
        sine[944] = -11'sd482;
        sine[945] = -11'sd476;
        sine[946] = -11'sd471;
        sine[947] = -11'sd465;
        sine[948] = -11'sd459;
        sine[949] = -11'sd454;
        sine[950] = -11'sd448;
        sine[951] = -11'sd443;
        sine[952] = -11'sd437;
        sine[953] = -11'sd431;
        sine[954] = -11'sd426;
        sine[955] = -11'sd420;
        sine[956] = -11'sd414;
        sine[957] = -11'sd408;
        sine[958] = -11'sd403;
        sine[959] = -11'sd397;
        sine[960] = -11'sd391;
        sine[961] = -11'sd385;
        sine[962] = -11'sd379;
        sine[963] = -11'sd374;
        sine[964] = -11'sd368;
        sine[965] = -11'sd362;
        sine[966] = -11'sd356;
        sine[967] = -11'sd350;
        sine[968] = -11'sd344;
        sine[969] = -11'sd338;
        sine[970] = -11'sd332;
        sine[971] = -11'sd326;
        sine[972] = -11'sd320;
        sine[973] = -11'sd314;
        sine[974] = -11'sd308;
        sine[975] = -11'sd302;
        sine[976] = -11'sd296;
        sine[977] = -11'sd290;
        sine[978] = -11'sd284;
        sine[979] = -11'sd278;
        sine[980] = -11'sd272;
        sine[981] = -11'sd266;
        sine[982] = -11'sd260;
        sine[983] = -11'sd254;
        sine[984] = -11'sd248;
        sine[985] = -11'sd242;
        sine[986] = -11'sd236;
        sine[987] = -11'sd230;
        sine[988] = -11'sd224;
        sine[989] = -11'sd218;
        sine[990] = -11'sd211;
        sine[991] = -11'sd205;
        sine[992] = -11'sd199;
        sine[993] = -11'sd193;
        sine[994] = -11'sd187;
        sine[995] = -11'sd181;
        sine[996] = -11'sd174;
        sine[997] = -11'sd168;
        sine[998] = -11'sd162;
        sine[999] = -11'sd156;
        sine[1000] = -11'sd150;
        sine[1001] = -11'sd143;
        sine[1002] = -11'sd137;
        sine[1003] = -11'sd131;
        sine[1004] = -11'sd125;
        sine[1005] = -11'sd118;
        sine[1006] = -11'sd112;
        sine[1007] = -11'sd106;
        sine[1008] = -11'sd100;
        sine[1009] = -11'sd94;
        sine[1010] = -11'sd87;
        sine[1011] = -11'sd81;
        sine[1012] = -11'sd75;
        sine[1013] = -11'sd68;
        sine[1014] = -11'sd62;
        sine[1015] = -11'sd56;
        sine[1016] = -11'sd50;
        sine[1017] = -11'sd43;
        sine[1018] = -11'sd37;
        sine[1019] = -11'sd31;
        sine[1020] = -11'sd25;
        sine[1021] = -11'sd18;
        sine[1022] = -11'sd12;
        sine[1023] = -11'sd6;
    end

endmodule


