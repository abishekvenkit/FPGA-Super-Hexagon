module tan(input  logic Clk,
           input  logic [9:0] angle,
           output logic [19:0] answer);

    reg signed [19:0] tangent [0:1023];

    always_ff @ (posedge Clk) begin
        answer <= tangent[angle];
    end

    initial begin
        tangent[0] = 20'sd0;
        tangent[1] = 20'sd6;
        tangent[2] = 20'sd12;
        tangent[3] = 20'sd18;
        tangent[4] = 20'sd25;
        tangent[5] = 20'sd31;
        tangent[6] = 20'sd37;
        tangent[7] = 20'sd44;
        tangent[8] = 20'sd50;
        tangent[9] = 20'sd56;
        tangent[10] = 20'sd62;
        tangent[11] = 20'sd69;
        tangent[12] = 20'sd75;
        tangent[13] = 20'sd81;
        tangent[14] = 20'sd88;
        tangent[15] = 20'sd94;
        tangent[16] = 20'sd100;
        tangent[17] = 20'sd107;
        tangent[18] = 20'sd113;
        tangent[19] = 20'sd119;
        tangent[20] = 20'sd126;
        tangent[21] = 20'sd132;
        tangent[22] = 20'sd139;
        tangent[23] = 20'sd145;
        tangent[24] = 20'sd151;
        tangent[25] = 20'sd158;
        tangent[26] = 20'sd164;
        tangent[27] = 20'sd171;
        tangent[28] = 20'sd177;
        tangent[29] = 20'sd184;
        tangent[30] = 20'sd190;
        tangent[31] = 20'sd197;
        tangent[32] = 20'sd203;
        tangent[33] = 20'sd210;
        tangent[34] = 20'sd216;
        tangent[35] = 20'sd223;
        tangent[36] = 20'sd229;
        tangent[37] = 20'sd236;
        tangent[38] = 20'sd243;
        tangent[39] = 20'sd249;
        tangent[40] = 20'sd256;
        tangent[41] = 20'sd263;
        tangent[42] = 20'sd269;
        tangent[43] = 20'sd276;
        tangent[44] = 20'sd283;
        tangent[45] = 20'sd290;
        tangent[46] = 20'sd296;
        tangent[47] = 20'sd303;
        tangent[48] = 20'sd310;
        tangent[49] = 20'sd317;
        tangent[50] = 20'sd324;
        tangent[51] = 20'sd331;
        tangent[52] = 20'sd338;
        tangent[53] = 20'sd345;
        tangent[54] = 20'sd352;
        tangent[55] = 20'sd359;
        tangent[56] = 20'sd366;
        tangent[57] = 20'sd373;
        tangent[58] = 20'sd380;
        tangent[59] = 20'sd387;
        tangent[60] = 20'sd395;
        tangent[61] = 20'sd402;
        tangent[62] = 20'sd409;
        tangent[63] = 20'sd416;
        tangent[64] = 20'sd424;
        tangent[65] = 20'sd431;
        tangent[66] = 20'sd438;
        tangent[67] = 20'sd446;
        tangent[68] = 20'sd453;
        tangent[69] = 20'sd461;
        tangent[70] = 20'sd469;
        tangent[71] = 20'sd476;
        tangent[72] = 20'sd484;
        tangent[73] = 20'sd492;
        tangent[74] = 20'sd499;
        tangent[75] = 20'sd507;
        tangent[76] = 20'sd515;
        tangent[77] = 20'sd523;
        tangent[78] = 20'sd531;
        tangent[79] = 20'sd539;
        tangent[80] = 20'sd547;
        tangent[81] = 20'sd555;
        tangent[82] = 20'sd563;
        tangent[83] = 20'sd571;
        tangent[84] = 20'sd580;
        tangent[85] = 20'sd588;
        tangent[86] = 20'sd596;
        tangent[87] = 20'sd605;
        tangent[88] = 20'sd613;
        tangent[89] = 20'sd622;
        tangent[90] = 20'sd630;
        tangent[91] = 20'sd639;
        tangent[92] = 20'sd648;
        tangent[93] = 20'sd657;
        tangent[94] = 20'sd666;
        tangent[95] = 20'sd675;
        tangent[96] = 20'sd684;
        tangent[97] = 20'sd693;
        tangent[98] = 20'sd702;
        tangent[99] = 20'sd711;
        tangent[100] = 20'sd721;
        tangent[101] = 20'sd730;
        tangent[102] = 20'sd740;
        tangent[103] = 20'sd749;
        tangent[104] = 20'sd759;
        tangent[105] = 20'sd769;
        tangent[106] = 20'sd779;
        tangent[107] = 20'sd789;
        tangent[108] = 20'sd799;
        tangent[109] = 20'sd809;
        tangent[110] = 20'sd819;
        tangent[111] = 20'sd829;
        tangent[112] = 20'sd840;
        tangent[113] = 20'sd850;
        tangent[114] = 20'sd861;
        tangent[115] = 20'sd872;
        tangent[116] = 20'sd883;
        tangent[117] = 20'sd894;
        tangent[118] = 20'sd905;
        tangent[119] = 20'sd916;
        tangent[120] = 20'sd928;
        tangent[121] = 20'sd939;
        tangent[122] = 20'sd951;
        tangent[123] = 20'sd963;
        tangent[124] = 20'sd974;
        tangent[125] = 20'sd986;
        tangent[126] = 20'sd999;
        tangent[127] = 20'sd1011;
        tangent[128] = 20'sd1023;
        tangent[129] = 20'sd1036;
        tangent[130] = 20'sd1049;
        tangent[131] = 20'sd1062;
        tangent[132] = 20'sd1075;
        tangent[133] = 20'sd1088;
        tangent[134] = 20'sd1102;
        tangent[135] = 20'sd1115;
        tangent[136] = 20'sd1129;
        tangent[137] = 20'sd1143;
        tangent[138] = 20'sd1158;
        tangent[139] = 20'sd1172;
        tangent[140] = 20'sd1187;
        tangent[141] = 20'sd1201;
        tangent[142] = 20'sd1216;
        tangent[143] = 20'sd1232;
        tangent[144] = 20'sd1247;
        tangent[145] = 20'sd1263;
        tangent[146] = 20'sd1279;
        tangent[147] = 20'sd1295;
        tangent[148] = 20'sd1312;
        tangent[149] = 20'sd1328;
        tangent[150] = 20'sd1345;
        tangent[151] = 20'sd1363;
        tangent[152] = 20'sd1380;
        tangent[153] = 20'sd1398;
        tangent[154] = 20'sd1416;
        tangent[155] = 20'sd1435;
        tangent[156] = 20'sd1453;
        tangent[157] = 20'sd1473;
        tangent[158] = 20'sd1492;
        tangent[159] = 20'sd1512;
        tangent[160] = 20'sd1532;
        tangent[161] = 20'sd1553;
        tangent[162] = 20'sd1574;
        tangent[163] = 20'sd1595;
        tangent[164] = 20'sd1617;
        tangent[165] = 20'sd1639;
        tangent[166] = 20'sd1661;
        tangent[167] = 20'sd1684;
        tangent[168] = 20'sd1708;
        tangent[169] = 20'sd1732;
        tangent[170] = 20'sd1756;
        tangent[171] = 20'sd1782;
        tangent[172] = 20'sd1807;
        tangent[173] = 20'sd1833;
        tangent[174] = 20'sd1860;
        tangent[175] = 20'sd1887;
        tangent[176] = 20'sd1915;
        tangent[177] = 20'sd1944;
        tangent[178] = 20'sd1973;
        tangent[179] = 20'sd2003;
        tangent[180] = 20'sd2034;
        tangent[181] = 20'sd2065;
        tangent[182] = 20'sd2098;
        tangent[183] = 20'sd2131;
        tangent[184] = 20'sd2165;
        tangent[185] = 20'sd2199;
        tangent[186] = 20'sd2235;
        tangent[187] = 20'sd2272;
        tangent[188] = 20'sd2310;
        tangent[189] = 20'sd2348;
        tangent[190] = 20'sd2388;
        tangent[191] = 20'sd2429;
        tangent[192] = 20'sd2472;
        tangent[193] = 20'sd2515;
        tangent[194] = 20'sd2560;
        tangent[195] = 20'sd2606;
        tangent[196] = 20'sd2654;
        tangent[197] = 20'sd2703;
        tangent[198] = 20'sd2754;
        tangent[199] = 20'sd2807;
        tangent[200] = 20'sd2861;
        tangent[201] = 20'sd2918;
        tangent[202] = 20'sd2976;
        tangent[203] = 20'sd3036;
        tangent[204] = 20'sd3099;
        tangent[205] = 20'sd3164;
        tangent[206] = 20'sd3232;
        tangent[207] = 20'sd3302;
        tangent[208] = 20'sd3375;
        tangent[209] = 20'sd3451;
        tangent[210] = 20'sd3531;
        tangent[211] = 20'sd3613;
        tangent[212] = 20'sd3700;
        tangent[213] = 20'sd3790;
        tangent[214] = 20'sd3885;
        tangent[215] = 20'sd3984;
        tangent[216] = 20'sd4088;
        tangent[217] = 20'sd4197;
        tangent[218] = 20'sd4311;
        tangent[219] = 20'sd4432;
        tangent[220] = 20'sd4560;
        tangent[221] = 20'sd4694;
        tangent[222] = 20'sd4836;
        tangent[223] = 20'sd4987;
        tangent[224] = 20'sd5147;
        tangent[225] = 20'sd5318;
        tangent[226] = 20'sd5499;
        tangent[227] = 20'sd5693;
        tangent[228] = 20'sd5901;
        tangent[229] = 20'sd6124;
        tangent[230] = 20'sd6364;
        tangent[231] = 20'sd6622;
        tangent[232] = 20'sd6903;
        tangent[233] = 20'sd7207;
        tangent[234] = 20'sd7539;
        tangent[235] = 20'sd7902;
        tangent[236] = 20'sd8302;
        tangent[237] = 20'sd8743;
        tangent[238] = 20'sd9233;
        tangent[239] = 20'sd9781;
        tangent[240] = 20'sd10396;
        tangent[241] = 20'sd11094;
        tangent[242] = 20'sd11891;
        tangent[243] = 20'sd12810;
        tangent[244] = 20'sd13882;
        tangent[245] = 20'sd15148;
        tangent[246] = 20'sd16667;
        tangent[247] = 20'sd18524;
        tangent[248] = 20'sd20843;
        tangent[249] = 20'sd23826;
        tangent[250] = 20'sd27801;
        tangent[251] = 20'sd33366;
        tangent[252] = 20'sd41713;
        tangent[253] = 20'sd55622;
        tangent[254] = 20'sd83438;
        tangent[255] = 20'sd166883;
        tangent[256] = 20'sd524287;
        tangent[257] = -20'sd166883;
        tangent[258] = -20'sd83438;
        tangent[259] = -20'sd55622;
        tangent[260] = -20'sd41713;
        tangent[261] = -20'sd33366;
        tangent[262] = -20'sd27801;
        tangent[263] = -20'sd23826;
        tangent[264] = -20'sd20843;
        tangent[265] = -20'sd18524;
        tangent[266] = -20'sd16667;
        tangent[267] = -20'sd15148;
        tangent[268] = -20'sd13882;
        tangent[269] = -20'sd12810;
        tangent[270] = -20'sd11891;
        tangent[271] = -20'sd11094;
        tangent[272] = -20'sd10396;
        tangent[273] = -20'sd9781;
        tangent[274] = -20'sd9233;
        tangent[275] = -20'sd8743;
        tangent[276] = -20'sd8302;
        tangent[277] = -20'sd7902;
        tangent[278] = -20'sd7539;
        tangent[279] = -20'sd7207;
        tangent[280] = -20'sd6903;
        tangent[281] = -20'sd6622;
        tangent[282] = -20'sd6364;
        tangent[283] = -20'sd6124;
        tangent[284] = -20'sd5901;
        tangent[285] = -20'sd5693;
        tangent[286] = -20'sd5499;
        tangent[287] = -20'sd5318;
        tangent[288] = -20'sd5147;
        tangent[289] = -20'sd4987;
        tangent[290] = -20'sd4836;
        tangent[291] = -20'sd4694;
        tangent[292] = -20'sd4560;
        tangent[293] = -20'sd4432;
        tangent[294] = -20'sd4311;
        tangent[295] = -20'sd4197;
        tangent[296] = -20'sd4088;
        tangent[297] = -20'sd3984;
        tangent[298] = -20'sd3885;
        tangent[299] = -20'sd3790;
        tangent[300] = -20'sd3700;
        tangent[301] = -20'sd3613;
        tangent[302] = -20'sd3531;
        tangent[303] = -20'sd3451;
        tangent[304] = -20'sd3375;
        tangent[305] = -20'sd3302;
        tangent[306] = -20'sd3232;
        tangent[307] = -20'sd3164;
        tangent[308] = -20'sd3099;
        tangent[309] = -20'sd3036;
        tangent[310] = -20'sd2976;
        tangent[311] = -20'sd2918;
        tangent[312] = -20'sd2861;
        tangent[313] = -20'sd2807;
        tangent[314] = -20'sd2754;
        tangent[315] = -20'sd2703;
        tangent[316] = -20'sd2654;
        tangent[317] = -20'sd2606;
        tangent[318] = -20'sd2560;
        tangent[319] = -20'sd2515;
        tangent[320] = -20'sd2472;
        tangent[321] = -20'sd2429;
        tangent[322] = -20'sd2388;
        tangent[323] = -20'sd2348;
        tangent[324] = -20'sd2310;
        tangent[325] = -20'sd2272;
        tangent[326] = -20'sd2235;
        tangent[327] = -20'sd2199;
        tangent[328] = -20'sd2165;
        tangent[329] = -20'sd2131;
        tangent[330] = -20'sd2098;
        tangent[331] = -20'sd2065;
        tangent[332] = -20'sd2034;
        tangent[333] = -20'sd2003;
        tangent[334] = -20'sd1973;
        tangent[335] = -20'sd1944;
        tangent[336] = -20'sd1915;
        tangent[337] = -20'sd1887;
        tangent[338] = -20'sd1860;
        tangent[339] = -20'sd1833;
        tangent[340] = -20'sd1807;
        tangent[341] = -20'sd1782;
        tangent[342] = -20'sd1756;
        tangent[343] = -20'sd1732;
        tangent[344] = -20'sd1708;
        tangent[345] = -20'sd1684;
        tangent[346] = -20'sd1661;
        tangent[347] = -20'sd1639;
        tangent[348] = -20'sd1617;
        tangent[349] = -20'sd1595;
        tangent[350] = -20'sd1574;
        tangent[351] = -20'sd1553;
        tangent[352] = -20'sd1532;
        tangent[353] = -20'sd1512;
        tangent[354] = -20'sd1492;
        tangent[355] = -20'sd1473;
        tangent[356] = -20'sd1453;
        tangent[357] = -20'sd1435;
        tangent[358] = -20'sd1416;
        tangent[359] = -20'sd1398;
        tangent[360] = -20'sd1380;
        tangent[361] = -20'sd1363;
        tangent[362] = -20'sd1345;
        tangent[363] = -20'sd1328;
        tangent[364] = -20'sd1312;
        tangent[365] = -20'sd1295;
        tangent[366] = -20'sd1279;
        tangent[367] = -20'sd1263;
        tangent[368] = -20'sd1247;
        tangent[369] = -20'sd1232;
        tangent[370] = -20'sd1216;
        tangent[371] = -20'sd1201;
        tangent[372] = -20'sd1187;
        tangent[373] = -20'sd1172;
        tangent[374] = -20'sd1158;
        tangent[375] = -20'sd1143;
        tangent[376] = -20'sd1129;
        tangent[377] = -20'sd1115;
        tangent[378] = -20'sd1102;
        tangent[379] = -20'sd1088;
        tangent[380] = -20'sd1075;
        tangent[381] = -20'sd1062;
        tangent[382] = -20'sd1049;
        tangent[383] = -20'sd1036;
        tangent[384] = -20'sd1024;
        tangent[385] = -20'sd1011;
        tangent[386] = -20'sd999;
        tangent[387] = -20'sd986;
        tangent[388] = -20'sd974;
        tangent[389] = -20'sd963;
        tangent[390] = -20'sd951;
        tangent[391] = -20'sd939;
        tangent[392] = -20'sd928;
        tangent[393] = -20'sd916;
        tangent[394] = -20'sd905;
        tangent[395] = -20'sd894;
        tangent[396] = -20'sd883;
        tangent[397] = -20'sd872;
        tangent[398] = -20'sd861;
        tangent[399] = -20'sd850;
        tangent[400] = -20'sd840;
        tangent[401] = -20'sd829;
        tangent[402] = -20'sd819;
        tangent[403] = -20'sd809;
        tangent[404] = -20'sd799;
        tangent[405] = -20'sd789;
        tangent[406] = -20'sd779;
        tangent[407] = -20'sd769;
        tangent[408] = -20'sd759;
        tangent[409] = -20'sd749;
        tangent[410] = -20'sd740;
        tangent[411] = -20'sd730;
        tangent[412] = -20'sd721;
        tangent[413] = -20'sd711;
        tangent[414] = -20'sd702;
        tangent[415] = -20'sd693;
        tangent[416] = -20'sd684;
        tangent[417] = -20'sd675;
        tangent[418] = -20'sd666;
        tangent[419] = -20'sd657;
        tangent[420] = -20'sd648;
        tangent[421] = -20'sd639;
        tangent[422] = -20'sd630;
        tangent[423] = -20'sd622;
        tangent[424] = -20'sd613;
        tangent[425] = -20'sd605;
        tangent[426] = -20'sd596;
        tangent[427] = -20'sd588;
        tangent[428] = -20'sd580;
        tangent[429] = -20'sd571;
        tangent[430] = -20'sd563;
        tangent[431] = -20'sd555;
        tangent[432] = -20'sd547;
        tangent[433] = -20'sd539;
        tangent[434] = -20'sd531;
        tangent[435] = -20'sd523;
        tangent[436] = -20'sd515;
        tangent[437] = -20'sd507;
        tangent[438] = -20'sd499;
        tangent[439] = -20'sd492;
        tangent[440] = -20'sd484;
        tangent[441] = -20'sd476;
        tangent[442] = -20'sd469;
        tangent[443] = -20'sd461;
        tangent[444] = -20'sd453;
        tangent[445] = -20'sd446;
        tangent[446] = -20'sd438;
        tangent[447] = -20'sd431;
        tangent[448] = -20'sd424;
        tangent[449] = -20'sd416;
        tangent[450] = -20'sd409;
        tangent[451] = -20'sd402;
        tangent[452] = -20'sd395;
        tangent[453] = -20'sd387;
        tangent[454] = -20'sd380;
        tangent[455] = -20'sd373;
        tangent[456] = -20'sd366;
        tangent[457] = -20'sd359;
        tangent[458] = -20'sd352;
        tangent[459] = -20'sd345;
        tangent[460] = -20'sd338;
        tangent[461] = -20'sd331;
        tangent[462] = -20'sd324;
        tangent[463] = -20'sd317;
        tangent[464] = -20'sd310;
        tangent[465] = -20'sd303;
        tangent[466] = -20'sd296;
        tangent[467] = -20'sd290;
        tangent[468] = -20'sd283;
        tangent[469] = -20'sd276;
        tangent[470] = -20'sd269;
        tangent[471] = -20'sd263;
        tangent[472] = -20'sd256;
        tangent[473] = -20'sd249;
        tangent[474] = -20'sd243;
        tangent[475] = -20'sd236;
        tangent[476] = -20'sd229;
        tangent[477] = -20'sd223;
        tangent[478] = -20'sd216;
        tangent[479] = -20'sd210;
        tangent[480] = -20'sd203;
        tangent[481] = -20'sd197;
        tangent[482] = -20'sd190;
        tangent[483] = -20'sd184;
        tangent[484] = -20'sd177;
        tangent[485] = -20'sd171;
        tangent[486] = -20'sd164;
        tangent[487] = -20'sd158;
        tangent[488] = -20'sd151;
        tangent[489] = -20'sd145;
        tangent[490] = -20'sd139;
        tangent[491] = -20'sd132;
        tangent[492] = -20'sd126;
        tangent[493] = -20'sd119;
        tangent[494] = -20'sd113;
        tangent[495] = -20'sd107;
        tangent[496] = -20'sd100;
        tangent[497] = -20'sd94;
        tangent[498] = -20'sd88;
        tangent[499] = -20'sd81;
        tangent[500] = -20'sd75;
        tangent[501] = -20'sd69;
        tangent[502] = -20'sd62;
        tangent[503] = -20'sd56;
        tangent[504] = -20'sd50;
        tangent[505] = -20'sd44;
        tangent[506] = -20'sd37;
        tangent[507] = -20'sd31;
        tangent[508] = -20'sd25;
        tangent[509] = -20'sd18;
        tangent[510] = -20'sd12;
        tangent[511] = -20'sd6;
        tangent[512] = 20'sd0;
        tangent[513] = 20'sd6;
        tangent[514] = 20'sd12;
        tangent[515] = 20'sd18;
        tangent[516] = 20'sd25;
        tangent[517] = 20'sd31;
        tangent[518] = 20'sd37;
        tangent[519] = 20'sd44;
        tangent[520] = 20'sd50;
        tangent[521] = 20'sd56;
        tangent[522] = 20'sd62;
        tangent[523] = 20'sd69;
        tangent[524] = 20'sd75;
        tangent[525] = 20'sd81;
        tangent[526] = 20'sd88;
        tangent[527] = 20'sd94;
        tangent[528] = 20'sd100;
        tangent[529] = 20'sd107;
        tangent[530] = 20'sd113;
        tangent[531] = 20'sd119;
        tangent[532] = 20'sd126;
        tangent[533] = 20'sd132;
        tangent[534] = 20'sd139;
        tangent[535] = 20'sd145;
        tangent[536] = 20'sd151;
        tangent[537] = 20'sd158;
        tangent[538] = 20'sd164;
        tangent[539] = 20'sd171;
        tangent[540] = 20'sd177;
        tangent[541] = 20'sd184;
        tangent[542] = 20'sd190;
        tangent[543] = 20'sd197;
        tangent[544] = 20'sd203;
        tangent[545] = 20'sd210;
        tangent[546] = 20'sd216;
        tangent[547] = 20'sd223;
        tangent[548] = 20'sd229;
        tangent[549] = 20'sd236;
        tangent[550] = 20'sd243;
        tangent[551] = 20'sd249;
        tangent[552] = 20'sd256;
        tangent[553] = 20'sd263;
        tangent[554] = 20'sd269;
        tangent[555] = 20'sd276;
        tangent[556] = 20'sd283;
        tangent[557] = 20'sd290;
        tangent[558] = 20'sd296;
        tangent[559] = 20'sd303;
        tangent[560] = 20'sd310;
        tangent[561] = 20'sd317;
        tangent[562] = 20'sd324;
        tangent[563] = 20'sd331;
        tangent[564] = 20'sd338;
        tangent[565] = 20'sd345;
        tangent[566] = 20'sd352;
        tangent[567] = 20'sd359;
        tangent[568] = 20'sd366;
        tangent[569] = 20'sd373;
        tangent[570] = 20'sd380;
        tangent[571] = 20'sd387;
        tangent[572] = 20'sd395;
        tangent[573] = 20'sd402;
        tangent[574] = 20'sd409;
        tangent[575] = 20'sd416;
        tangent[576] = 20'sd424;
        tangent[577] = 20'sd431;
        tangent[578] = 20'sd438;
        tangent[579] = 20'sd446;
        tangent[580] = 20'sd453;
        tangent[581] = 20'sd461;
        tangent[582] = 20'sd469;
        tangent[583] = 20'sd476;
        tangent[584] = 20'sd484;
        tangent[585] = 20'sd492;
        tangent[586] = 20'sd499;
        tangent[587] = 20'sd507;
        tangent[588] = 20'sd515;
        tangent[589] = 20'sd523;
        tangent[590] = 20'sd531;
        tangent[591] = 20'sd539;
        tangent[592] = 20'sd547;
        tangent[593] = 20'sd555;
        tangent[594] = 20'sd563;
        tangent[595] = 20'sd571;
        tangent[596] = 20'sd580;
        tangent[597] = 20'sd588;
        tangent[598] = 20'sd596;
        tangent[599] = 20'sd605;
        tangent[600] = 20'sd613;
        tangent[601] = 20'sd622;
        tangent[602] = 20'sd630;
        tangent[603] = 20'sd639;
        tangent[604] = 20'sd648;
        tangent[605] = 20'sd657;
        tangent[606] = 20'sd666;
        tangent[607] = 20'sd675;
        tangent[608] = 20'sd684;
        tangent[609] = 20'sd693;
        tangent[610] = 20'sd702;
        tangent[611] = 20'sd711;
        tangent[612] = 20'sd721;
        tangent[613] = 20'sd730;
        tangent[614] = 20'sd740;
        tangent[615] = 20'sd749;
        tangent[616] = 20'sd759;
        tangent[617] = 20'sd769;
        tangent[618] = 20'sd779;
        tangent[619] = 20'sd789;
        tangent[620] = 20'sd799;
        tangent[621] = 20'sd809;
        tangent[622] = 20'sd819;
        tangent[623] = 20'sd829;
        tangent[624] = 20'sd840;
        tangent[625] = 20'sd850;
        tangent[626] = 20'sd861;
        tangent[627] = 20'sd872;
        tangent[628] = 20'sd883;
        tangent[629] = 20'sd894;
        tangent[630] = 20'sd905;
        tangent[631] = 20'sd916;
        tangent[632] = 20'sd928;
        tangent[633] = 20'sd939;
        tangent[634] = 20'sd951;
        tangent[635] = 20'sd963;
        tangent[636] = 20'sd974;
        tangent[637] = 20'sd986;
        tangent[638] = 20'sd999;
        tangent[639] = 20'sd1011;
        tangent[640] = 20'sd1023;
        tangent[641] = 20'sd1036;
        tangent[642] = 20'sd1049;
        tangent[643] = 20'sd1062;
        tangent[644] = 20'sd1075;
        tangent[645] = 20'sd1088;
        tangent[646] = 20'sd1102;
        tangent[647] = 20'sd1115;
        tangent[648] = 20'sd1129;
        tangent[649] = 20'sd1143;
        tangent[650] = 20'sd1158;
        tangent[651] = 20'sd1172;
        tangent[652] = 20'sd1187;
        tangent[653] = 20'sd1201;
        tangent[654] = 20'sd1216;
        tangent[655] = 20'sd1232;
        tangent[656] = 20'sd1247;
        tangent[657] = 20'sd1263;
        tangent[658] = 20'sd1279;
        tangent[659] = 20'sd1295;
        tangent[660] = 20'sd1312;
        tangent[661] = 20'sd1328;
        tangent[662] = 20'sd1345;
        tangent[663] = 20'sd1363;
        tangent[664] = 20'sd1380;
        tangent[665] = 20'sd1398;
        tangent[666] = 20'sd1416;
        tangent[667] = 20'sd1435;
        tangent[668] = 20'sd1453;
        tangent[669] = 20'sd1473;
        tangent[670] = 20'sd1492;
        tangent[671] = 20'sd1512;
        tangent[672] = 20'sd1532;
        tangent[673] = 20'sd1553;
        tangent[674] = 20'sd1574;
        tangent[675] = 20'sd1595;
        tangent[676] = 20'sd1617;
        tangent[677] = 20'sd1639;
        tangent[678] = 20'sd1661;
        tangent[679] = 20'sd1684;
        tangent[680] = 20'sd1708;
        tangent[681] = 20'sd1732;
        tangent[682] = 20'sd1756;
        tangent[683] = 20'sd1782;
        tangent[684] = 20'sd1807;
        tangent[685] = 20'sd1833;
        tangent[686] = 20'sd1860;
        tangent[687] = 20'sd1887;
        tangent[688] = 20'sd1915;
        tangent[689] = 20'sd1944;
        tangent[690] = 20'sd1973;
        tangent[691] = 20'sd2003;
        tangent[692] = 20'sd2034;
        tangent[693] = 20'sd2065;
        tangent[694] = 20'sd2098;
        tangent[695] = 20'sd2131;
        tangent[696] = 20'sd2165;
        tangent[697] = 20'sd2199;
        tangent[698] = 20'sd2235;
        tangent[699] = 20'sd2272;
        tangent[700] = 20'sd2310;
        tangent[701] = 20'sd2348;
        tangent[702] = 20'sd2388;
        tangent[703] = 20'sd2429;
        tangent[704] = 20'sd2472;
        tangent[705] = 20'sd2515;
        tangent[706] = 20'sd2560;
        tangent[707] = 20'sd2606;
        tangent[708] = 20'sd2654;
        tangent[709] = 20'sd2703;
        tangent[710] = 20'sd2754;
        tangent[711] = 20'sd2807;
        tangent[712] = 20'sd2861;
        tangent[713] = 20'sd2918;
        tangent[714] = 20'sd2976;
        tangent[715] = 20'sd3036;
        tangent[716] = 20'sd3099;
        tangent[717] = 20'sd3164;
        tangent[718] = 20'sd3232;
        tangent[719] = 20'sd3302;
        tangent[720] = 20'sd3375;
        tangent[721] = 20'sd3451;
        tangent[722] = 20'sd3531;
        tangent[723] = 20'sd3613;
        tangent[724] = 20'sd3700;
        tangent[725] = 20'sd3790;
        tangent[726] = 20'sd3885;
        tangent[727] = 20'sd3984;
        tangent[728] = 20'sd4088;
        tangent[729] = 20'sd4197;
        tangent[730] = 20'sd4311;
        tangent[731] = 20'sd4432;
        tangent[732] = 20'sd4560;
        tangent[733] = 20'sd4694;
        tangent[734] = 20'sd4836;
        tangent[735] = 20'sd4987;
        tangent[736] = 20'sd5147;
        tangent[737] = 20'sd5318;
        tangent[738] = 20'sd5499;
        tangent[739] = 20'sd5693;
        tangent[740] = 20'sd5901;
        tangent[741] = 20'sd6124;
        tangent[742] = 20'sd6364;
        tangent[743] = 20'sd6622;
        tangent[744] = 20'sd6903;
        tangent[745] = 20'sd7207;
        tangent[746] = 20'sd7539;
        tangent[747] = 20'sd7902;
        tangent[748] = 20'sd8302;
        tangent[749] = 20'sd8743;
        tangent[750] = 20'sd9233;
        tangent[751] = 20'sd9781;
        tangent[752] = 20'sd10396;
        tangent[753] = 20'sd11094;
        tangent[754] = 20'sd11891;
        tangent[755] = 20'sd12810;
        tangent[756] = 20'sd13882;
        tangent[757] = 20'sd15148;
        tangent[758] = 20'sd16667;
        tangent[759] = 20'sd18524;
        tangent[760] = 20'sd20843;
        tangent[761] = 20'sd23826;
        tangent[762] = 20'sd27801;
        tangent[763] = 20'sd33366;
        tangent[764] = 20'sd41713;
        tangent[765] = 20'sd55622;
        tangent[766] = 20'sd83438;
        tangent[767] = 20'sd166883;
        tangent[768] = 20'sd524287;
        tangent[769] = -20'sd166883;
        tangent[770] = -20'sd83438;
        tangent[771] = -20'sd55622;
        tangent[772] = -20'sd41713;
        tangent[773] = -20'sd33366;
        tangent[774] = -20'sd27801;
        tangent[775] = -20'sd23826;
        tangent[776] = -20'sd20843;
        tangent[777] = -20'sd18524;
        tangent[778] = -20'sd16667;
        tangent[779] = -20'sd15148;
        tangent[780] = -20'sd13882;
        tangent[781] = -20'sd12810;
        tangent[782] = -20'sd11891;
        tangent[783] = -20'sd11094;
        tangent[784] = -20'sd10396;
        tangent[785] = -20'sd9781;
        tangent[786] = -20'sd9233;
        tangent[787] = -20'sd8743;
        tangent[788] = -20'sd8302;
        tangent[789] = -20'sd7902;
        tangent[790] = -20'sd7539;
        tangent[791] = -20'sd7207;
        tangent[792] = -20'sd6903;
        tangent[793] = -20'sd6622;
        tangent[794] = -20'sd6364;
        tangent[795] = -20'sd6124;
        tangent[796] = -20'sd5901;
        tangent[797] = -20'sd5693;
        tangent[798] = -20'sd5499;
        tangent[799] = -20'sd5318;
        tangent[800] = -20'sd5147;
        tangent[801] = -20'sd4987;
        tangent[802] = -20'sd4836;
        tangent[803] = -20'sd4694;
        tangent[804] = -20'sd4560;
        tangent[805] = -20'sd4432;
        tangent[806] = -20'sd4311;
        tangent[807] = -20'sd4197;
        tangent[808] = -20'sd4088;
        tangent[809] = -20'sd3984;
        tangent[810] = -20'sd3885;
        tangent[811] = -20'sd3790;
        tangent[812] = -20'sd3700;
        tangent[813] = -20'sd3613;
        tangent[814] = -20'sd3531;
        tangent[815] = -20'sd3451;
        tangent[816] = -20'sd3375;
        tangent[817] = -20'sd3302;
        tangent[818] = -20'sd3232;
        tangent[819] = -20'sd3164;
        tangent[820] = -20'sd3099;
        tangent[821] = -20'sd3036;
        tangent[822] = -20'sd2976;
        tangent[823] = -20'sd2918;
        tangent[824] = -20'sd2861;
        tangent[825] = -20'sd2807;
        tangent[826] = -20'sd2754;
        tangent[827] = -20'sd2703;
        tangent[828] = -20'sd2654;
        tangent[829] = -20'sd2606;
        tangent[830] = -20'sd2560;
        tangent[831] = -20'sd2515;
        tangent[832] = -20'sd2472;
        tangent[833] = -20'sd2429;
        tangent[834] = -20'sd2388;
        tangent[835] = -20'sd2348;
        tangent[836] = -20'sd2310;
        tangent[837] = -20'sd2272;
        tangent[838] = -20'sd2235;
        tangent[839] = -20'sd2199;
        tangent[840] = -20'sd2165;
        tangent[841] = -20'sd2131;
        tangent[842] = -20'sd2098;
        tangent[843] = -20'sd2065;
        tangent[844] = -20'sd2034;
        tangent[845] = -20'sd2003;
        tangent[846] = -20'sd1973;
        tangent[847] = -20'sd1944;
        tangent[848] = -20'sd1915;
        tangent[849] = -20'sd1887;
        tangent[850] = -20'sd1860;
        tangent[851] = -20'sd1833;
        tangent[852] = -20'sd1807;
        tangent[853] = -20'sd1782;
        tangent[854] = -20'sd1756;
        tangent[855] = -20'sd1732;
        tangent[856] = -20'sd1708;
        tangent[857] = -20'sd1684;
        tangent[858] = -20'sd1661;
        tangent[859] = -20'sd1639;
        tangent[860] = -20'sd1617;
        tangent[861] = -20'sd1595;
        tangent[862] = -20'sd1574;
        tangent[863] = -20'sd1553;
        tangent[864] = -20'sd1532;
        tangent[865] = -20'sd1512;
        tangent[866] = -20'sd1492;
        tangent[867] = -20'sd1473;
        tangent[868] = -20'sd1453;
        tangent[869] = -20'sd1435;
        tangent[870] = -20'sd1416;
        tangent[871] = -20'sd1398;
        tangent[872] = -20'sd1380;
        tangent[873] = -20'sd1363;
        tangent[874] = -20'sd1345;
        tangent[875] = -20'sd1328;
        tangent[876] = -20'sd1312;
        tangent[877] = -20'sd1295;
        tangent[878] = -20'sd1279;
        tangent[879] = -20'sd1263;
        tangent[880] = -20'sd1247;
        tangent[881] = -20'sd1232;
        tangent[882] = -20'sd1216;
        tangent[883] = -20'sd1201;
        tangent[884] = -20'sd1187;
        tangent[885] = -20'sd1172;
        tangent[886] = -20'sd1158;
        tangent[887] = -20'sd1143;
        tangent[888] = -20'sd1129;
        tangent[889] = -20'sd1115;
        tangent[890] = -20'sd1102;
        tangent[891] = -20'sd1088;
        tangent[892] = -20'sd1075;
        tangent[893] = -20'sd1062;
        tangent[894] = -20'sd1049;
        tangent[895] = -20'sd1036;
        tangent[896] = -20'sd1024;
        tangent[897] = -20'sd1011;
        tangent[898] = -20'sd999;
        tangent[899] = -20'sd986;
        tangent[900] = -20'sd974;
        tangent[901] = -20'sd963;
        tangent[902] = -20'sd951;
        tangent[903] = -20'sd939;
        tangent[904] = -20'sd928;
        tangent[905] = -20'sd916;
        tangent[906] = -20'sd905;
        tangent[907] = -20'sd894;
        tangent[908] = -20'sd883;
        tangent[909] = -20'sd872;
        tangent[910] = -20'sd861;
        tangent[911] = -20'sd850;
        tangent[912] = -20'sd840;
        tangent[913] = -20'sd829;
        tangent[914] = -20'sd819;
        tangent[915] = -20'sd809;
        tangent[916] = -20'sd799;
        tangent[917] = -20'sd789;
        tangent[918] = -20'sd779;
        tangent[919] = -20'sd769;
        tangent[920] = -20'sd759;
        tangent[921] = -20'sd749;
        tangent[922] = -20'sd740;
        tangent[923] = -20'sd730;
        tangent[924] = -20'sd721;
        tangent[925] = -20'sd711;
        tangent[926] = -20'sd702;
        tangent[927] = -20'sd693;
        tangent[928] = -20'sd684;
        tangent[929] = -20'sd675;
        tangent[930] = -20'sd666;
        tangent[931] = -20'sd657;
        tangent[932] = -20'sd648;
        tangent[933] = -20'sd639;
        tangent[934] = -20'sd630;
        tangent[935] = -20'sd622;
        tangent[936] = -20'sd613;
        tangent[937] = -20'sd605;
        tangent[938] = -20'sd596;
        tangent[939] = -20'sd588;
        tangent[940] = -20'sd580;
        tangent[941] = -20'sd571;
        tangent[942] = -20'sd563;
        tangent[943] = -20'sd555;
        tangent[944] = -20'sd547;
        tangent[945] = -20'sd539;
        tangent[946] = -20'sd531;
        tangent[947] = -20'sd523;
        tangent[948] = -20'sd515;
        tangent[949] = -20'sd507;
        tangent[950] = -20'sd499;
        tangent[951] = -20'sd492;
        tangent[952] = -20'sd484;
        tangent[953] = -20'sd476;
        tangent[954] = -20'sd469;
        tangent[955] = -20'sd461;
        tangent[956] = -20'sd453;
        tangent[957] = -20'sd446;
        tangent[958] = -20'sd438;
        tangent[959] = -20'sd431;
        tangent[960] = -20'sd424;
        tangent[961] = -20'sd416;
        tangent[962] = -20'sd409;
        tangent[963] = -20'sd402;
        tangent[964] = -20'sd395;
        tangent[965] = -20'sd387;
        tangent[966] = -20'sd380;
        tangent[967] = -20'sd373;
        tangent[968] = -20'sd366;
        tangent[969] = -20'sd359;
        tangent[970] = -20'sd352;
        tangent[971] = -20'sd345;
        tangent[972] = -20'sd338;
        tangent[973] = -20'sd331;
        tangent[974] = -20'sd324;
        tangent[975] = -20'sd317;
        tangent[976] = -20'sd310;
        tangent[977] = -20'sd303;
        tangent[978] = -20'sd296;
        tangent[979] = -20'sd290;
        tangent[980] = -20'sd283;
        tangent[981] = -20'sd276;
        tangent[982] = -20'sd269;
        tangent[983] = -20'sd263;
        tangent[984] = -20'sd256;
        tangent[985] = -20'sd249;
        tangent[986] = -20'sd243;
        tangent[987] = -20'sd236;
        tangent[988] = -20'sd229;
        tangent[989] = -20'sd223;
        tangent[990] = -20'sd216;
        tangent[991] = -20'sd210;
        tangent[992] = -20'sd203;
        tangent[993] = -20'sd197;
        tangent[994] = -20'sd190;
        tangent[995] = -20'sd184;
        tangent[996] = -20'sd177;
        tangent[997] = -20'sd171;
        tangent[998] = -20'sd164;
        tangent[999] = -20'sd158;
        tangent[1000] = -20'sd151;
        tangent[1001] = -20'sd145;
        tangent[1002] = -20'sd139;
        tangent[1003] = -20'sd132;
        tangent[1004] = -20'sd126;
        tangent[1005] = -20'sd119;
        tangent[1006] = -20'sd113;
        tangent[1007] = -20'sd107;
        tangent[1008] = -20'sd100;
        tangent[1009] = -20'sd94;
        tangent[1010] = -20'sd88;
        tangent[1011] = -20'sd81;
        tangent[1012] = -20'sd75;
        tangent[1013] = -20'sd69;
        tangent[1014] = -20'sd62;
        tangent[1015] = -20'sd56;
        tangent[1016] = -20'sd50;
        tangent[1017] = -20'sd44;
        tangent[1018] = -20'sd37;
        tangent[1019] = -20'sd31;
        tangent[1020] = -20'sd25;
        tangent[1021] = -20'sd18;
        tangent[1022] = -20'sd12;
        tangent[1023] = -20'sd6;
    end

endmodule